// This is a generated file. Use and modify at your own risk.
//////////////////////////////////////////////////////////////////////////////// 
// default_nettype of none prevents implicit wire declaration.
`include "accelerator.vh"
`default_nettype none
module delta_pr_accelerator_axi_top #(
  parameter integer C_M00_AXI_ADDR_WIDTH = 64 ,
  parameter integer C_M00_AXI_DATA_WIDTH = 512,
  parameter integer C_M01_AXI_ADDR_WIDTH = 64 ,
  parameter integer C_M01_AXI_DATA_WIDTH = 512,
  // acc parameter
  parameter integer V_ID_WIDTH = `V_ID_WIDTH,
  parameter integer V_OFF_AWIDTH = `V_OFF_AWIDTH,
  parameter integer V_OFF_DWIDTH = `V_OFF_DWIDTH,
  parameter integer V_VALUE_WIDTH = `V_VALUE_WIDTH,
  parameter integer CORE_NUM = `CORE_NUM,
  parameter integer CORE_NUM_WIDTH = `CORE_NUM_WIDTH,
  parameter integer ITERATION_WIDTH = `ITERATION_WIDTH,
  parameter integer HBM_AWIDTH = `HBM_AWIDTH,
  parameter integer HBM_DWIDTH = `HBM_DWIDTH,
  parameter integer HBM_DWIDTH_PER_CORE = `HBM_DWIDTH_PER_CORE,
  parameter integer HBM_EDGE_MASK = `HBM_EDGE_MASK,
  parameter integer PSEUDO_CHANNEL_NUM = `PSEUDO_CHANNEL_NUM,
  parameter integer GROUP_CORE_NUM = `GROUP_CORE_NUM,
  parameter integer DELTA_BRAM_AWIDTH = `DELTA_BRAM_AWIDTH
)
(
  // System Signals
  input  wire                              ap_clk         ,
  input  wire                              ap_rst_n       ,
  // AXI4 master interface m00_axi
  output wire                              m00_axi_awvalid,
  input  wire                              m00_axi_awready,
  output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_awaddr ,
  output wire [8-1:0]                      m00_axi_awlen  ,
  output wire                              m00_axi_wvalid ,
  input  wire                              m00_axi_wready ,
  output wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_wdata  ,
  output wire [C_M00_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb  ,
  output wire                              m00_axi_wlast  ,
  input  wire                              m00_axi_bvalid ,
  output wire                              m00_axi_bready ,
  output wire                              m00_axi_arvalid,
  input  wire                              m00_axi_arready,
  output wire [C_M00_AXI_ADDR_WIDTH-1:0]   m00_axi_araddr ,
  output wire [8-1:0]                      m00_axi_arlen  ,
  input  wire                              m00_axi_rvalid ,
  output wire                              m00_axi_rready ,
  input  wire [C_M00_AXI_DATA_WIDTH-1:0]   m00_axi_rdata  ,
  input  wire                              m00_axi_rlast  ,
  // AXI4 master interface m01_axi
  output wire                              m01_axi_awvalid,
  input  wire                              m01_axi_awready,
  output wire [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_awaddr ,
  output wire [8-1:0]                      m01_axi_awlen  ,
  output wire                              m01_axi_wvalid ,
  input  wire                              m01_axi_wready ,
  output wire [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_wdata  ,
  output wire [C_M01_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb  ,
  output wire                              m01_axi_wlast  ,
  input  wire                              m01_axi_bvalid ,
  output wire                              m01_axi_bready ,
  output wire                              m01_axi_arvalid,
  input  wire                              m01_axi_arready,
  output wire [C_M01_AXI_ADDR_WIDTH-1:0]   m01_axi_araddr ,
  output wire [8-1:0]                      m01_axi_arlen  ,
  input  wire                              m01_axi_rvalid ,
  output wire                              m01_axi_rready ,
  input  wire [C_M01_AXI_DATA_WIDTH-1:0]   m01_axi_rdata  ,
  input  wire                              m01_axi_rlast  ,
  // Control Signals
  input  wire                              ap_start       ,
  output wire                              ap_idle        ,
  output wire                              ap_done        ,
  output wire                              ap_ready       ,
  input  wire [32-1:0]                     one_over_n     ,
  input  wire [32-1:0]                     added_const    ,
  input  wire [32-1:0]                     delta2_value   ,//reg????????????????//
  input  wire [32-1:0]                     bitmap_compressed_num,
  input  wire [64-1:0]                     axi00_ptr0     ,
  input  wire [64-1:0]                     axi01_ptr0     
);


timeunit 1ps;
timeprecision 1ps;

///////////////////////////////////////////////////////////////////////////////
// Local Parameters
///////////////////////////////////////////////////////////////////////////////
// Large enough for interesting traffic.
localparam integer  LP_DEFAULT_LENGTH_IN_BYTES = 16384;
localparam integer  LP_NUM_EXAMPLES    = 2;

///////////////////////////////////////////////////////////////////////////////
// Wires and Variables
///////////////////////////////////////////////////////////////////////////////
(* KEEP = "yes" *)
logic                                areset                         = 1'b0;
logic                                ap_start_r                     = 1'b0;
logic                                ap_idle_r                      = 1'b1;
logic                                ap_start_pulse                ;
logic [LP_NUM_EXAMPLES-1:0]          ap_done_i                     ;
logic [LP_NUM_EXAMPLES-1:0]          ap_done_r                      = {LP_NUM_EXAMPLES{1'b0}};
logic [32-1:0]                       ctrl_constant                  = 32'd1;
// kernel
wire [CORE_NUM - 1 : 0]                 P1_iteration_done;
wire [CORE_NUM - 1 : 0]                 P1_next_rst;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P1_active_v_id;
wire [CORE_NUM - 1 : 0]                 P1_active_v_valid;
wire [CORE_NUM - 1 : 0]                 P1_iteration_end;
wire [CORE_NUM - 1 : 0]                 P1_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0]  P1_iteration_id;

wire [CORE_NUM - 1 : 0]                 P2_next_rst;
wire [CORE_NUM - 1 : 0]                 P2_stage_full;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P2_active_v_id;
wire [CORE_NUM - 1 : 0]                 P2_active_v_id_valid;
wire [CORE_NUM * V_OFF_AWIDTH - 1 : 0]  P2_rd_active_v_offset_addr;
wire [CORE_NUM * DELTA_BRAM_AWIDTH - 1 : 0]  P2_rd_active_v_value_addr;
wire [CORE_NUM - 1 : 0]                 P2_rd_active_v_addr_valid;
wire [CORE_NUM - 1 : 0]                 P2_iteration_end;
wire [CORE_NUM - 1 : 0]                 P2_iteration_end_valid;
wire [CORE_NUM *ITERATION_WIDTH - 1 : 0]P2_iteration_id;

wire [CORE_NUM - 1 : 0]                 P3_transfer_complete;
wire [PSEUDO_CHANNEL_NUM * HBM_AWIDTH - 1 : 0]  P3_hbm_controller_addr;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]  P3_hbm_addr_valid;
wire [CORE_NUM - 1 : 0]                 P3_next_rst;
wire [CORE_NUM * V_OFF_DWIDTH - 1 : 0]  P3_active_v_loffset;
wire [CORE_NUM * V_OFF_DWIDTH - 1 : 0]  P3_active_v_roffset;
wire [CORE_NUM - 1 : 0]                 P3_active_v_valid;

wire [CORE_NUM - 1 : 0]                 P4_next_rst;
wire [CORE_NUM - 1 : 0]                 P4_stage_full;
wire [CORE_NUM * HBM_AWIDTH - 1 : 0]    P4_rd_hbm_edge_addr;
wire [CORE_NUM * HBM_EDGE_MASK - 1 : 0] P4_rd_hbm_edge_mask;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P4_hbm_active_v_id;
wire [CORE_NUM - 1 : 0]                 P4_rd_hbm_edge_valid;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0] P4_hbm_active_v_value;
wire [CORE_NUM - 1 : 0]                 P4_hbm_active_v_value_valid;
wire [CORE_NUM - 1 : 0]                 P4_iteration_end;
wire [CORE_NUM - 1 : 0]                 P4_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0]  P4_iteration_id;

wire [CORE_NUM - 1 : 0]                 P5_next_rst;
wire [CORE_NUM - 1 : 0]                 P5_stage_full;
wire [PSEUDO_CHANNEL_NUM * HBM_AWIDTH - 1 : 0]    P5_rd_hbm_edge_addr;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]                 P5_rd_hbm_edge_valid;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P5_active_v_id;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0] P5_active_v_value;
wire [CORE_NUM - 1 : 0]                 P5_active_v_valid;
wire [CORE_NUM - 1 : 0]                 P5_iteration_end;
wire [CORE_NUM - 1 : 0]                 P5_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0]  P5_iteration_id;

wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_interface_full;
wire [PSEUDO_CHANNEL_NUM * HBM_AWIDTH - 1 : 0]  HBM_interface_rd_hbm_edge_addr;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_interface_rd_hbm_edge_valid;
wire [CORE_NUM * HBM_AWIDTH - 1 : 0]  HBM_interface_active_v_edge;
wire [CORE_NUM - 1 : 0]               HBM_interface_active_v_edge_valid;

wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_controller_read_full;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_controller_write_full;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_controller_write_empty;
wire [PSEUDO_CHANNEL_NUM * HBM_DWIDTH - 1 : 0]  HBM_controller_edge;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_controller_valid;
wire [PSEUDO_CHANNEL_NUM * HBM_AWIDTH - 1 : 0]  HBM_controller_recv_addr;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]               HBM_controller_addr_valid;

wire [CORE_NUM - 1 : 0]                 P7_next_rst;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]       P7_stage_full;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P7_update_v_id;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0] P7_update_v_value;
wire [CORE_NUM - 1 : 0]                 P7_update_v_valid;
wire [CORE_NUM - 1 : 0]                 P7_iteration_end;
wire [CORE_NUM - 1 : 0]                 P7_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0]  P7_iteration_id;

wire [CORE_NUM - 1 : 0]                 P8_next_rst;
wire [CORE_NUM - 1 : 0]                 P8_stage_full;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]    P8_update_v_id;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0] P8_update_v_value;
wire [CORE_NUM - 1 : 0]                 P8_update_v_valid;
wire [CORE_NUM - 1 : 0]                 P8_iteration_end;
wire [CORE_NUM - 1 : 0]                 P8_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0]  P8_iteration_id;

wire [CORE_NUM - 1 : 0]                   P9_next_rst;
wire [CORE_NUM - 1 : 0]                   P9_dest_core_full;
wire [CORE_NUM * V_OFF_AWIDTH - 1 : 0]      P9_wr_vertex_bram_addr;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0]   P9_wr_vertex_bram_data;
wire [CORE_NUM - 1 : 0]                   P9_wr_vertex_bram_valid;
wire [CORE_NUM - 1 : 0]                   P9_wr_vertex_bram_iteration_end;
wire [CORE_NUM - 1 : 0]                   P9_wr_vertex_bram_iteration_end_valid;
wire [CORE_NUM * ITERATION_WIDTH - 1 : 0] P9_wr_vertex_bram_iteration_id;

wire [CORE_NUM - 1 : 0]                   P10_next_rst;
wire                                      P10_transfer_done;
wire [CORE_NUM * HBM_DWIDTH_PER_CORE - 1 : 0] P10_wb_bfs_data;
wire [PSEUDO_CHANNEL_NUM - 1 : 0]             P10_wb_bfs_valid;
wire [CORE_NUM - 1 : 0]                   P10_stage_full;
wire [CORE_NUM * V_VALUE_WIDTH - 1 : 0]   P10_src_recv_update_v_value;
wire [CORE_NUM - 1 : 0]                   P10_src_recv_update_v_valid;
wire [CORE_NUM * V_ID_WIDTH - 1 : 0]      P10_backend_active_v_id;
wire [CORE_NUM - 1 : 0]                   P10_backend_active_v_updated;
wire [CORE_NUM - 1 : 0]                   P10_backend_active_v_valid;
wire [CORE_NUM - 1 : 0]                   P10_iteration_end;
wire [CORE_NUM - 1 : 0]                   P10_iteration_end_valid;

wire [CORE_NUM * V_ID_WIDTH - 1 : 0]      P11_active_v_id;
wire [CORE_NUM - 1 : 0]                   P11_active_v_updated;
wire [CORE_NUM - 1 : 0]                   P11_active_v_valid;
wire [CORE_NUM - 1 : 0]                   P11_iteration_end;
wire [CORE_NUM - 1 : 0]                   P11_iteration_end_valid;

// 8 vertex per channel, 64bit per vertex : 32 for value, 32 for id
wire [32 * 16 - 1 : 0] WR_BACK_bfs_res [0 : LP_NUM_EXAMPLES - 1];
wire WR_BACK_bfs_valid [0 : LP_NUM_EXAMPLES - 1];

(* keep = "TRUE" *)   wire          clk = ap_clk;
reg rst, uram_rst, cycle_valid;
reg [31 : 0] acc_cycle;
reg [2 : 0] acc_state; // 00: initial state; 01: transfer uram data; 10: running; 11: done
wire transfer_uram;
wire transfer_bram;
assign transfer_uram = (acc_state == 2'b01);
assign transfer_bram = (acc_state == 2'b11); // transfer bram data after acc done

always @ (posedge clk) begin
  if (areset) begin
    acc_state <= 2'b00;
    rst <= 1'b1;
    uram_rst <= 1'b1;
  end else begin
    case (acc_state)
      2'b00: if (ap_start_pulse) begin
        acc_state <= 2'b01;
        rst <= 1'b1;
        uram_rst <= 1'b0;
      end
      2'b01: if (P3_transfer_complete == {CORE_NUM{1'b1}}) begin
        acc_state <= 2'b10;
        rst <= 1'b0;
        uram_rst <= 1'b0;
      end
      2'b10: if (P1_iteration_done == {CORE_NUM{1'b1}}) begin
        acc_state <= 2'b11;
        rst <= 1'b1;
        uram_rst <= 1'b0;
      end
      2'b11: begin
        // keep done signal
      end
    endcase
  end
end

// BUFG u_AXI_CLK_IN_0  ( .I (ap_clk), .O (clk) );

///////////////////////////////////////////////////////////////////////////////
// Begin RTL
///////////////////////////////////////////////////////////////////////////////

//cycle inc
always @(posedge ap_clk) begin
  if(acc_state < 2) begin
    acc_cycle <= 0;
  end else if (acc_state == 2) begin
    acc_cycle <= acc_cycle + 1;
  end
  if(acc_state < 3 && P1_iteration_done != {CORE_NUM{1'b1}}) begin
    cycle_valid <=0;
  end else if(acc_state == 2 && P1_iteration_done == {CORE_NUM{1'b1}}) begin
    cycle_valid <=1;
  end else if (acc_state == 3) begin
    cycle_valid <=0;
  end
end

// Register and invert reset signal.
always @(posedge ap_clk) begin
  areset <= ~ap_rst_n;
end

// create pulse when ap_start transitions to 1
always @(posedge ap_clk) begin
  begin
    ap_start_r <= ap_start;
  end
end

assign ap_start_pulse = ap_start & ~ap_start_r;

// ap_idle is asserted when done is asserted, it is de-asserted when ap_start_pulse
// is asserted
always @(posedge ap_clk) begin
  if (areset) begin
    ap_idle_r <= 1'b1;
  end
  else begin
    ap_idle_r <= ap_done ? 1'b1 :
      ap_start_pulse ? 1'b0 : ap_idle;
  end
end

assign ap_idle = ap_idle_r;

// Done logic
always @(posedge ap_clk) begin
  if (areset) begin
    ap_done_r <= '0;
  end
  else begin
    ap_done_r <= (ap_done) ? '0 : ap_done_r | ap_done_i;
  end
end

assign ap_done = &ap_done_r && (acc_state == 2'b11) && P10_transfer_done;

// Ready Logic (non-pipelined case)
assign ap_ready = ap_done;

// combine result
generate
  genvar i;
  for (i = 0; i < PSEUDO_CHANNEL_NUM; i = i + 1) begin
    assign WR_BACK_bfs_res[i] = P10_wb_bfs_data[(i + 1) * HBM_DWIDTH - 1 : i * HBM_DWIDTH];
    assign WR_BACK_bfs_valid[i] = P10_wb_bfs_valid[i];
  end
endgenerate

assign HBM_controller_recv_addr = transfer_uram ? P3_hbm_controller_addr : HBM_interface_rd_hbm_edge_addr;
assign HBM_controller_addr_valid = transfer_uram ? P3_hbm_addr_valid : HBM_interface_rd_hbm_edge_valid;

// HBM controller
hbm_channel_controller #(
  .C_M_AXI_ADDR_WIDTH ( C_M00_AXI_ADDR_WIDTH ),
  .C_M_AXI_DATA_WIDTH ( C_M00_AXI_DATA_WIDTH ),
  .C_ADDER_BIT_WIDTH  ( 32                   )
)
hbm_channel_controller_inst_m00_axi (
  .aclk                    ( ap_clk                  ),
  .areset                  ( areset                  ),
  .kernel_clk              ( ap_clk                  ),
  .kernel_rst              ( areset                  ),
  .ctrl_addr_offset        ( axi00_ptr0              ),
  .ctrl_constant           ( ctrl_constant           ),
  .ap_start                ( ap_start_pulse          ),
  .m_axi_awvalid           ( m00_axi_awvalid         ),
  .m_axi_awready           ( m00_axi_awready         ),
  .m_axi_awaddr            ( m00_axi_awaddr          ),
  .m_axi_awlen             ( m00_axi_awlen           ),
  .m_axi_wvalid            ( m00_axi_wvalid          ),
  .m_axi_wready            ( m00_axi_wready          ),
  .m_axi_wdata             ( m00_axi_wdata           ),
  .m_axi_wstrb             ( m00_axi_wstrb           ),
  .m_axi_wlast             ( m00_axi_wlast           ),
  .m_axi_bvalid            ( m00_axi_bvalid          ),
  .m_axi_bready            ( m00_axi_bready          ),
  .m_axi_arvalid           ( m00_axi_arvalid         ),
  .m_axi_arready           ( m00_axi_arready         ),
  .m_axi_araddr            ( m00_axi_araddr          ),
  .m_axi_arlen             ( m00_axi_arlen           ),
  .m_axi_rvalid            ( m00_axi_rvalid          ),
  .m_axi_rready            ( m00_axi_rready          ),
  .m_axi_rdata             ( m00_axi_rdata           ),
  .m_axi_rlast             ( m00_axi_rlast           ),
  // acc
  .controller_recv_edge_addr        ({{32{1'b0}},HBM_controller_recv_addr[(0 + 1) * HBM_AWIDTH - 1 : 0 * HBM_AWIDTH]}<<6),
  .controller_recv_edge_addr_valid  (HBM_controller_addr_valid[0]),
  .read_stage_full                  (HBM_controller_read_full[0]),
  .controller_send_edge             (HBM_controller_edge[(0 + 1) * HBM_DWIDTH - 1 : 0 * HBM_DWIDTH]),
  .controller_send_edge_valid       (HBM_controller_valid[0]),
  .controller_recv_update_data      (cycle_valid ? {{480{1'b0}},acc_cycle} : WR_BACK_bfs_res[0]),
  .controller_recv_update_addr      (), // not use, should increment internal
  .controller_recv_update_valid     (cycle_valid ? 1'b1 : |WR_BACK_bfs_valid[0]),
  .write_stage_full                 (HBM_controller_write_full[0]),
  .write_stage_empty                (ap_done_i[0])
);

hbm_channel_controller #(
  .C_M_AXI_ADDR_WIDTH ( C_M01_AXI_ADDR_WIDTH ),
  .C_M_AXI_DATA_WIDTH ( C_M01_AXI_DATA_WIDTH ),
  .C_ADDER_BIT_WIDTH  ( 32                   )
)
hbm_channel_controller_inst_m01_axi (
  .aclk                    ( ap_clk                  ),
  .areset                  ( areset                  ),
  .kernel_clk              ( ap_clk                  ),
  .kernel_rst              ( areset                  ),
  .ctrl_addr_offset        ( axi01_ptr0              ),
  .ctrl_constant           ( ctrl_constant           ),
  .ap_start                ( ap_start_pulse          ),
  .m_axi_awvalid           ( m01_axi_awvalid         ),
  .m_axi_awready           ( m01_axi_awready         ),
  .m_axi_awaddr            ( m01_axi_awaddr          ),
  .m_axi_awlen             ( m01_axi_awlen           ),
  .m_axi_wvalid            ( m01_axi_wvalid          ),
  .m_axi_wready            ( m01_axi_wready          ),
  .m_axi_wdata             ( m01_axi_wdata           ),
  .m_axi_wstrb             ( m01_axi_wstrb           ),
  .m_axi_wlast             ( m01_axi_wlast           ),
  .m_axi_bvalid            ( m01_axi_bvalid          ),
  .m_axi_bready            ( m01_axi_bready          ),
  .m_axi_arvalid           ( m01_axi_arvalid         ),
  .m_axi_arready           ( m01_axi_arready         ),
  .m_axi_araddr            ( m01_axi_araddr          ),
  .m_axi_arlen             ( m01_axi_arlen           ),
  .m_axi_rvalid            ( m01_axi_rvalid          ),
  .m_axi_rready            ( m01_axi_rready          ),
  .m_axi_rdata             ( m01_axi_rdata           ),
  .m_axi_rlast             ( m01_axi_rlast           ),
  // acc
  .controller_recv_edge_addr        ({{32{1'b0}},HBM_controller_recv_addr[(1 + 1) * HBM_AWIDTH - 1 : 1 * HBM_AWIDTH]}<<6),
  .controller_recv_edge_addr_valid  (HBM_controller_addr_valid[1]),
  .read_stage_full                  (HBM_controller_read_full[1]),
  .controller_send_edge             (HBM_controller_edge[(1 + 1) * HBM_DWIDTH - 1 : 1 * HBM_DWIDTH]),
  .controller_send_edge_valid       (HBM_controller_valid[1]),
  .controller_recv_update_data      (WR_BACK_bfs_res[1]),
  .controller_recv_update_addr      (), // not use, should increment internal
  .controller_recv_update_valid     (|WR_BACK_bfs_valid[1]),
  .write_stage_full                 (HBM_controller_write_full[1]),
  .write_stage_empty                (ap_done_i[1])
);


// kernel
rd_active_vertex  RD_ACTIVE_VERTEX (
  .clk                (clk),
  .rst                (rst),
  .bitmap_compressed_num      (bitmap_compressed_num),
  .backend_active_v_id        (P11_active_v_id),
  .backend_active_v_updated   (P11_active_v_updated),
  .backend_active_v_id_valid  (P11_active_v_valid),
  .backend_iteration_end      (P11_iteration_end),
  .backend_iteration_end_valid(P11_iteration_end_valid),
  .next_stage_full            (P2_stage_full),

  .next_rst                   (P1_next_rst),
  .iteration_done             (P1_iteration_done),
  .active_v_id                (P1_active_v_id),
  .active_v_id_valid          (P1_active_v_valid),
  .iteration_end              (P1_iteration_end),
  .iteration_end_valid        (P1_iteration_end_valid),
  .iteration_id               (P1_iteration_id)
);

rd_active_vertex_offset RD_ACTIVE_VERTEX_OFFSET (
  .clk                        (clk),
  .rst                        (P1_next_rst),
  .front_active_v_id          (P1_active_v_id),
  .front_active_v_valid       (P1_active_v_valid),
  .front_iteration_end        (P1_iteration_end),
  .front_iteration_end_valid  (P1_iteration_end_valid),
  .front_iteration_id         (P1_iteration_id),
  .next_stage_full            (P4_stage_full),

  .next_rst                   (P2_next_rst),
  .stage_full                 (P2_stage_full),
  .active_v_id                (P2_active_v_id),
  .active_v_id_valid          (P2_active_v_id_valid),
  .rd_active_v_offset_addr    (P2_rd_active_v_offset_addr),
  .rd_active_v_value_addr     (P2_rd_active_v_value_addr),
  .rd_active_v_addr_valid     (P2_rd_active_v_addr_valid),
  .iteration_end              (P2_iteration_end),
  .iteration_end_valid        (P2_iteration_end_valid),
  .iteration_id               (P2_iteration_id)
);

offset_uram OFFSET_URAM (
  .clk                        (clk),
  .uram_rst                   (uram_rst),
  .hbm_controller_data        (HBM_controller_edge),
  .hbm_data_valid             (transfer_uram ? HBM_controller_valid : 0),
  .hbm_controller_full        (HBM_controller_read_full),
  .rst                        (P2_next_rst),
  .front_rd_active_v_offset_addr  (P2_rd_active_v_offset_addr),
  .front_active_v_valid       (P2_rd_active_v_addr_valid),

  .hbm_controller_addr        (P3_hbm_controller_addr),
  .hbm_addr_valid             (P3_hbm_addr_valid),
  .transfer_complete          (P3_transfer_complete),
  .next_rst                   (P3_next_rst),
  .uram_loffset               (P3_active_v_loffset),
  .uram_roffset               (P3_active_v_roffset),
  .uram_dvalid                (P3_active_v_valid)
);

rd_active_vertex_edge RD_ACTIVE_VERTEX_EDGE (
  .clk                        (clk),
  .rst                        (P2_next_rst),
  .front_active_v_id          (P2_active_v_id),
  .front_active_v_valid       (P2_active_v_id_valid),
  .front_active_v_loffset     (P3_active_v_loffset),
  .front_active_v_roffset     (P3_active_v_roffset),
  .front_offset_valid         (P3_active_v_valid),
  .front_iteration_end        (P2_iteration_end),
  .front_iteration_end_valid  (P2_iteration_end_valid),
  .front_iteration_id         (P2_iteration_id),
  .front_active_v_value       (P10_src_recv_update_v_value),
  .front_active_v_value_valid (P10_src_recv_update_v_valid),
  .combine_stage_full         (P5_stage_full),

  .next_rst                   (P4_next_rst),
  .stage_full                 (P4_stage_full),
  .rd_hbm_edge_addr           (P4_rd_hbm_edge_addr),
  .rd_hbm_edge_mask           (P4_rd_hbm_edge_mask),
  .hbm_active_v_id            (P4_hbm_active_v_id),
  .rd_hbm_edge_valid          (P4_rd_hbm_edge_valid),
  .hbm_active_v_value         (P4_hbm_active_v_value),
  .hbm_active_v_value_valid   (P4_hbm_active_v_value_valid),
  .iteration_end              (P4_iteration_end),
  .iteration_end_valid        (P4_iteration_end_valid),
  .iteration_id               (P4_iteration_id)
);

generate_hbm_edge_rqst GENERATE_HBM_EDGE_RQST (
  .clk                        (clk),
  .rst                        (P4_next_rst),
  .front_rd_hbm_edge_addr     (P4_rd_hbm_edge_addr),
  .front_rd_hbm_edge_mask     (P4_rd_hbm_edge_mask),
  .front_active_v_id          (P4_hbm_active_v_id),
  .front_rd_hbm_edge_valid    (P4_rd_hbm_edge_valid),
  .front_active_v_value       (P4_hbm_active_v_value),
  .front_active_v_value_valid (P4_hbm_active_v_value_valid),
  .front_iteration_end        (P4_iteration_end),
  .front_iteration_end_valid  (P4_iteration_end_valid),
  .front_iteration_id         (P4_iteration_id),
  .hbm_full                   (HBM_interface_full),
  .next_stage_full            (P7_stage_full),

  .next_rst                   (P5_next_rst),
  .stage_full                 (P5_stage_full),
  .rd_hbm_edge_addr           (P5_rd_hbm_edge_addr),
  .rd_hbm_edge_valid          (P5_rd_hbm_edge_valid),
  .active_v_id                (P5_active_v_id),
  .active_v_value             (P5_active_v_value),
  .active_v_id_valid          (P5_active_v_valid),
  .iteration_end              (P5_iteration_end),
  .iteration_end_valid        (P5_iteration_end_valid),
  .iteration_id               (P5_iteration_id)
);

hbm_interface HBM_INTERFACE (
  .clk                        (clk),
  .rst                        (P5_next_rst),
  .front_rd_hbm_edge_addr     (P5_rd_hbm_edge_addr),
  .front_rd_hbm_edge_valid    (P5_rd_hbm_edge_valid),
  .hbm_controller_edge        (HBM_controller_edge),
  .hbm_controller_valid       (HBM_controller_valid),
  .hbm_controller_full        (HBM_controller_read_full),

  .stage_full                 (HBM_interface_full),
  .rd_hbm_edge_addr           (HBM_interface_rd_hbm_edge_addr),
  .rd_hbm_edge_valid          (HBM_interface_rd_hbm_edge_valid),
  .active_v_edge              (HBM_interface_active_v_edge),
  .active_v_edge_valid        (HBM_interface_active_v_edge_valid)
);

scheduler SCHEDULER (
  .clk                        (clk),
  .rst                        (P5_next_rst),
  .front_active_v_id          (P5_active_v_id),
  .front_active_v_value       (P5_active_v_value),
  .front_active_v_valid       (P5_active_v_valid),
  .front_iteration_end        (P5_iteration_end),
  .front_iteration_end_valid  (P5_iteration_end_valid),
  .front_iteration_id         (P5_iteration_id),
  .hbm_interface_active_v_edge  (HBM_interface_active_v_edge),
  .hbm_interface_active_v_edge_valid  (HBM_interface_active_v_edge_valid),
  .next_stage_full            (P8_stage_full),

  .next_rst                   (P7_next_rst),
  .stage_full                 (P7_stage_full),
  .update_v_id                (P7_update_v_id),
  .update_v_value             (P7_update_v_value),
  .update_v_valid             (P7_update_v_valid),
  .iteration_end              (P7_iteration_end),
  .iteration_end_valid        (P7_iteration_end_valid),
  .iteration_id               (P7_iteration_id)
);

HyperX_Network HYPERX_NETWORK(
    .clk                     (clk),
    .hy1_front_rst           (P7_next_rst),
    .hy1_front_push_flag     ({CORE_NUM{1'b1}}),
    .hy1_front_update_v_id   (P7_update_v_id),
    .hy1_front_update_v_value          (P7_update_v_value),
    .hy1_front_pull_first_flag         (0),
    .hy1_front_update_v_valid          (P7_update_v_valid),
    .hy1_front_iteration_end           (P7_iteration_end),
    .hy1_front_iteration_end_valid     (P7_iteration_end_valid),
    .hy1_front_iteration_id            (P7_iteration_id),

    .hy2_front_rst                        (0),
    .hy2_front_push_flag                  (0),
    .hy2_front_update_v_id                (0),
    .hy2_front_update_v_value             (0),
    .hy2_front_pull_first_flag            (0),
    .hy2_front_update_v_valid             (0),
    .hy2_front_iteration_end              (0),
    .hy2_front_iteration_end_valid        (0),
    .source_core_full                     (P9_dest_core_full),

    .hy1_rst                              (P8_next_rst),
    .hy2_rst                              (),
    .hy1_stage_full                       (P8_stage_full),
    .hy2_stage_full                       (),

    .hy1_push_flag                       (),
    .hy1_update_v_id                       (P8_update_v_id),
    .hy1_update_v_value                       (P8_update_v_value),
    .hy1_pull_first_flag                       (),
    .hy1_update_v_valid                       (P8_update_v_valid),
    .hy1_iteration_end                       (P8_iteration_end),
    .hy1_iteration_end_valid                       (P8_iteration_end_valid),
    .hy1_iteration_id                       (P8_iteration_id),

    .hy2_push_flag                            (),
    .hy2_update_v_id                            (),
    .hy2_update_v_value                            (),
    .hy2_pull_first_flag                            (),
    .hy2_update_v_valid                            (),
    .hy2_iteration_end                            (),
    .hy2_iteration_end_valid                            ()
);


backend_core BACKEND_CORE (
  .clk                      (clk),
  .rst                      (P8_next_rst),
  .recv_update_v_id         (P8_update_v_id),
  .recv_update_v_value      (P8_update_v_value),
  .recv_update_v_valid      (P8_update_v_valid),
  .recv_iteration_end       (P8_iteration_end),
  .recv_iteration_end_valid (P8_iteration_end_valid),
  .recv_iteration_id        (P8_iteration_id),
  .next_stage_full          (P10_stage_full),

  .next_rst                 (P9_next_rst),
  .dest_core_full           (P9_dest_core_full),
  .wr_vertex_bram_addr      (P9_wr_vertex_bram_addr),
  .wr_vertex_bram_data      (P9_wr_vertex_bram_data),
  .wr_vertex_bram_valid     (P9_wr_vertex_bram_valid),
  .wr_vertex_bram_iteration_end       (P9_wr_vertex_bram_iteration_end),
  .wr_vertex_bram_iteration_end_valid (P9_wr_vertex_bram_iteration_end_valid),
  .wr_vertex_bram_iteration_id        (P9_wr_vertex_bram_iteration_id)
);

vtx_ram_controller VTX_RAM_CONTROLLER (
  .clk                        (clk),
  .added_const                (added_const),
  .one_over_n                 (one_over_n),
  .delta2_value               (delta2_value),
  .bitmap_compressed_num      (bitmap_compressed_num),
  .rst                        (transfer_bram ? {CORE_NUM{1'b0}} : P9_next_rst),
  .acc_state                  (acc_state),
  .transfer_bram              (transfer_bram),
  .initial_bram               (transfer_uram),
  .uram_rst                   (uram_rst),
  .hbm_write_full             (HBM_controller_write_full),
  .rd_addr_src                (P2_rd_active_v_value_addr),
  .rd_valid_src               (P2_rd_active_v_addr_valid),
  .wr_addr_dst                (P9_wr_vertex_bram_addr),
  .wr_v_value_dst             (P9_wr_vertex_bram_data),
  .wr_valid_dst               (P9_wr_vertex_bram_valid),
  .front_iteration_end        (P9_wr_vertex_bram_iteration_end),
  .front_iteration_end_valid  (P9_wr_vertex_bram_iteration_end_valid),
  .front_iteration_id         (P9_wr_vertex_bram_iteration_id),
  
  .next_rst                   (P10_next_rst),
  .transfer_done              (P10_transfer_done),
  .wb_bfs_data                (P10_wb_bfs_data),
  .wb_bfs_valid               (P10_wb_bfs_valid),

  .stage_full                 (P10_stage_full),
  .src_recv_update_v_value    (P10_src_recv_update_v_value),
  .src_recv_update_v_valid    (P10_src_recv_update_v_valid),
  .backend_active_v_id        (P10_backend_active_v_id),
  .backend_active_v_updated   (P10_backend_active_v_updated),
  .backend_active_v_valid     (P10_backend_active_v_valid),
  .iteration_end              (P10_iteration_end),
  .iteration_end_valid        (P10_iteration_end_valid)
);

apply_iteration_end APPLY_ITERATION_END (
  .clk                        (clk),
  .rst                        (P10_next_rst),
  .front_active_v_id          (P10_backend_active_v_id),
  .front_active_v_updated     (P10_backend_active_v_updated),
  .front_active_v_valid       (P10_backend_active_v_valid),
  .front_iteration_end        (P10_iteration_end),
  .front_iteration_end_valid  (P10_iteration_end_valid),

  .active_v_id                (P11_active_v_id),
  .active_v_updated           (P11_active_v_updated),
  .active_v_valid             (P11_active_v_valid),
  .iteration_end              (P11_iteration_end),
  .iteration_end_valid        (P11_iteration_end_valid)
);

endmodule : delta_pr_accelerator_axi_top
`default_nettype wire