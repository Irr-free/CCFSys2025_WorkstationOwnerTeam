// This is a generated file. Use and modify at your own risk.
////////////////////////////////////////////////////////////////////////////////
// default_nettype of none prevents implicit wire declaration.
`default_nettype none
`timescale 1 ps / 1 ps
import axi_vip_pkg::*;
import slv_m00_axi_vip_pkg::*;
import slv_m01_axi_vip_pkg::*;
import slv_m02_axi_vip_pkg::*;
import slv_m03_axi_vip_pkg::*;
import slv_m04_axi_vip_pkg::*;
import slv_m05_axi_vip_pkg::*;
import slv_m06_axi_vip_pkg::*;
import slv_m07_axi_vip_pkg::*;
import slv_m08_axi_vip_pkg::*;
import slv_m09_axi_vip_pkg::*;
import slv_m10_axi_vip_pkg::*;
import slv_m11_axi_vip_pkg::*;
import slv_m12_axi_vip_pkg::*;
import slv_m13_axi_vip_pkg::*;
import slv_m14_axi_vip_pkg::*;
import slv_m15_axi_vip_pkg::*;
import slv_m16_axi_vip_pkg::*;
import slv_m17_axi_vip_pkg::*;
import slv_m18_axi_vip_pkg::*;
import slv_m19_axi_vip_pkg::*;
import slv_m20_axi_vip_pkg::*;
import slv_m21_axi_vip_pkg::*;
import slv_m22_axi_vip_pkg::*;
import slv_m23_axi_vip_pkg::*;
import slv_m24_axi_vip_pkg::*;
import slv_m25_axi_vip_pkg::*;
import slv_m26_axi_vip_pkg::*;
import slv_m27_axi_vip_pkg::*;
import slv_m28_axi_vip_pkg::*;
import slv_m29_axi_vip_pkg::*;
import slv_m30_axi_vip_pkg::*;
import slv_m31_axi_vip_pkg::*;
import control_acc_kernel_vip_pkg::*;
module acc_kernel_tb ();
parameter integer LP_MAX_LENGTH = 8192;
parameter integer LP_MAX_TRANSFER_LENGTH = 16384 / 4;
parameter integer C_S_AXI_CONTROL_ADDR_WIDTH = 12;
parameter integer C_S_AXI_CONTROL_DATA_WIDTH = 32;
parameter integer C_M00_AXI_ADDR_WIDTH = 64;
parameter integer C_M00_AXI_DATA_WIDTH = 512;
parameter integer C_M01_AXI_ADDR_WIDTH = 64;
parameter integer C_M01_AXI_DATA_WIDTH = 512;
parameter integer C_M02_AXI_ADDR_WIDTH = 64;
parameter integer C_M02_AXI_DATA_WIDTH = 512;
parameter integer C_M03_AXI_ADDR_WIDTH = 64;
parameter integer C_M03_AXI_DATA_WIDTH = 512;
parameter integer C_M04_AXI_ADDR_WIDTH = 64;
parameter integer C_M04_AXI_DATA_WIDTH = 512;
parameter integer C_M05_AXI_ADDR_WIDTH = 64;
parameter integer C_M05_AXI_DATA_WIDTH = 512;
parameter integer C_M06_AXI_ADDR_WIDTH = 64;
parameter integer C_M06_AXI_DATA_WIDTH = 512;
parameter integer C_M07_AXI_ADDR_WIDTH = 64;
parameter integer C_M07_AXI_DATA_WIDTH = 512;
parameter integer C_M08_AXI_ADDR_WIDTH = 64;
parameter integer C_M08_AXI_DATA_WIDTH = 512;
parameter integer C_M09_AXI_ADDR_WIDTH = 64;
parameter integer C_M09_AXI_DATA_WIDTH = 512;
parameter integer C_M10_AXI_ADDR_WIDTH = 64;
parameter integer C_M10_AXI_DATA_WIDTH = 512;
parameter integer C_M11_AXI_ADDR_WIDTH = 64;
parameter integer C_M11_AXI_DATA_WIDTH = 512;
parameter integer C_M12_AXI_ADDR_WIDTH = 64;
parameter integer C_M12_AXI_DATA_WIDTH = 512;
parameter integer C_M13_AXI_ADDR_WIDTH = 64;
parameter integer C_M13_AXI_DATA_WIDTH = 512;
parameter integer C_M14_AXI_ADDR_WIDTH = 64;
parameter integer C_M14_AXI_DATA_WIDTH = 512;
parameter integer C_M15_AXI_ADDR_WIDTH = 64;
parameter integer C_M15_AXI_DATA_WIDTH = 512;
parameter integer C_M16_AXI_ADDR_WIDTH = 64;
parameter integer C_M16_AXI_DATA_WIDTH = 512;
parameter integer C_M17_AXI_ADDR_WIDTH = 64;
parameter integer C_M17_AXI_DATA_WIDTH = 512;
parameter integer C_M18_AXI_ADDR_WIDTH = 64;
parameter integer C_M18_AXI_DATA_WIDTH = 512;
parameter integer C_M19_AXI_ADDR_WIDTH = 64;
parameter integer C_M19_AXI_DATA_WIDTH = 512;
parameter integer C_M20_AXI_ADDR_WIDTH = 64;
parameter integer C_M20_AXI_DATA_WIDTH = 512;
parameter integer C_M21_AXI_ADDR_WIDTH = 64;
parameter integer C_M21_AXI_DATA_WIDTH = 512;
parameter integer C_M22_AXI_ADDR_WIDTH = 64;
parameter integer C_M22_AXI_DATA_WIDTH = 512;
parameter integer C_M23_AXI_ADDR_WIDTH = 64;
parameter integer C_M23_AXI_DATA_WIDTH = 512;
parameter integer C_M24_AXI_ADDR_WIDTH = 64;
parameter integer C_M24_AXI_DATA_WIDTH = 512;
parameter integer C_M25_AXI_ADDR_WIDTH = 64;
parameter integer C_M25_AXI_DATA_WIDTH = 512;
parameter integer C_M26_AXI_ADDR_WIDTH = 64;
parameter integer C_M26_AXI_DATA_WIDTH = 512;
parameter integer C_M27_AXI_ADDR_WIDTH = 64;
parameter integer C_M27_AXI_DATA_WIDTH = 512;
parameter integer C_M28_AXI_ADDR_WIDTH = 64;
parameter integer C_M28_AXI_DATA_WIDTH = 512;
parameter integer C_M29_AXI_ADDR_WIDTH = 64;
parameter integer C_M29_AXI_DATA_WIDTH = 512;
parameter integer C_M30_AXI_ADDR_WIDTH = 64;
parameter integer C_M30_AXI_DATA_WIDTH = 512;
parameter integer C_M31_AXI_ADDR_WIDTH = 64;
parameter integer C_M31_AXI_DATA_WIDTH = 512;

// Control Register
parameter KRNL_CTRL_REG_ADDR     = 32'h00000000;
parameter CTRL_START_MASK        = 32'h00000001;
parameter CTRL_DONE_MASK         = 32'h00000002;
parameter CTRL_IDLE_MASK         = 32'h00000004;
parameter CTRL_READY_MASK        = 32'h00000008;
parameter CTRL_CONTINUE_MASK     = 32'h00000010; // Only ap_ctrl_chain
parameter CTRL_AUTO_RESTART_MASK = 32'h00000080; // Not used

// Global Interrupt Enable Register
parameter KRNL_GIE_REG_ADDR      = 32'h00000004;
parameter GIE_GIE_MASK           = 32'h00000001;
// IP Interrupt Enable Register
parameter KRNL_IER_REG_ADDR      = 32'h00000008;
parameter IER_DONE_MASK          = 32'h00000001;
parameter IER_READY_MASK         = 32'h00000002;
// IP Interrupt Status Register
parameter KRNL_ISR_REG_ADDR      = 32'h0000000c;
parameter ISR_DONE_MASK          = 32'h00000001;
parameter ISR_READY_MASK         = 32'h00000002;

parameter integer LP_CLK_PERIOD_PS = 4000; // 250 MHz

//System Signals
logic ap_clk = 0;

initial begin: AP_CLK
  forever begin
    ap_clk = #(LP_CLK_PERIOD_PS/2) ~ap_clk;
  end
end
 
//System Signals
logic ap_rst_n = 0;
logic initial_reset  =0;

task automatic ap_rst_n_sequence(input integer unsigned width = 20);
  @(posedge ap_clk);
  #1ps;
  ap_rst_n = 0;
  repeat (width) @(posedge ap_clk);
  #1ps;
  ap_rst_n = 1;
endtask

initial begin: AP_RST
  ap_rst_n_sequence(50);
  initial_reset =1;
end
//AXI4 master interface m00_axi
wire [1-1:0] m00_axi_awvalid;
wire [1-1:0] m00_axi_awready;
wire [C_M00_AXI_ADDR_WIDTH-1:0] m00_axi_awaddr;
wire [8-1:0] m00_axi_awlen;
wire [1-1:0] m00_axi_wvalid;
wire [1-1:0] m00_axi_wready;
wire [C_M00_AXI_DATA_WIDTH-1:0] m00_axi_wdata;
wire [C_M00_AXI_DATA_WIDTH/8-1:0] m00_axi_wstrb;
wire [1-1:0] m00_axi_wlast;
wire [1-1:0] m00_axi_bvalid;
wire [1-1:0] m00_axi_bready;
wire [1-1:0] m00_axi_arvalid;
wire [1-1:0] m00_axi_arready;
wire [C_M00_AXI_ADDR_WIDTH-1:0] m00_axi_araddr;
wire [8-1:0] m00_axi_arlen;
wire [1-1:0] m00_axi_rvalid;
wire [1-1:0] m00_axi_rready;
wire [C_M00_AXI_DATA_WIDTH-1:0] m00_axi_rdata;
wire [1-1:0] m00_axi_rlast;
//AXI4 master interface m01_axi
wire [1-1:0] m01_axi_awvalid;
wire [1-1:0] m01_axi_awready;
wire [C_M01_AXI_ADDR_WIDTH-1:0] m01_axi_awaddr;
wire [8-1:0] m01_axi_awlen;
wire [1-1:0] m01_axi_wvalid;
wire [1-1:0] m01_axi_wready;
wire [C_M01_AXI_DATA_WIDTH-1:0] m01_axi_wdata;
wire [C_M01_AXI_DATA_WIDTH/8-1:0] m01_axi_wstrb;
wire [1-1:0] m01_axi_wlast;
wire [1-1:0] m01_axi_bvalid;
wire [1-1:0] m01_axi_bready;
wire [1-1:0] m01_axi_arvalid;
wire [1-1:0] m01_axi_arready;
wire [C_M01_AXI_ADDR_WIDTH-1:0] m01_axi_araddr;
wire [8-1:0] m01_axi_arlen;
wire [1-1:0] m01_axi_rvalid;
wire [1-1:0] m01_axi_rready;
wire [C_M01_AXI_DATA_WIDTH-1:0] m01_axi_rdata;
wire [1-1:0] m01_axi_rlast;
//AXI4 master interface m02_axi
wire [1-1:0] m02_axi_awvalid;
wire [1-1:0] m02_axi_awready;
wire [C_M02_AXI_ADDR_WIDTH-1:0] m02_axi_awaddr;
wire [8-1:0] m02_axi_awlen;
wire [1-1:0] m02_axi_wvalid;
wire [1-1:0] m02_axi_wready;
wire [C_M02_AXI_DATA_WIDTH-1:0] m02_axi_wdata;
wire [C_M02_AXI_DATA_WIDTH/8-1:0] m02_axi_wstrb;
wire [1-1:0] m02_axi_wlast;
wire [1-1:0] m02_axi_bvalid;
wire [1-1:0] m02_axi_bready;
wire [1-1:0] m02_axi_arvalid;
wire [1-1:0] m02_axi_arready;
wire [C_M02_AXI_ADDR_WIDTH-1:0] m02_axi_araddr;
wire [8-1:0] m02_axi_arlen;
wire [1-1:0] m02_axi_rvalid;
wire [1-1:0] m02_axi_rready;
wire [C_M02_AXI_DATA_WIDTH-1:0] m02_axi_rdata;
wire [1-1:0] m02_axi_rlast;
//AXI4 master interface m03_axi
wire [1-1:0] m03_axi_awvalid;
wire [1-1:0] m03_axi_awready;
wire [C_M03_AXI_ADDR_WIDTH-1:0] m03_axi_awaddr;
wire [8-1:0] m03_axi_awlen;
wire [1-1:0] m03_axi_wvalid;
wire [1-1:0] m03_axi_wready;
wire [C_M03_AXI_DATA_WIDTH-1:0] m03_axi_wdata;
wire [C_M03_AXI_DATA_WIDTH/8-1:0] m03_axi_wstrb;
wire [1-1:0] m03_axi_wlast;
wire [1-1:0] m03_axi_bvalid;
wire [1-1:0] m03_axi_bready;
wire [1-1:0] m03_axi_arvalid;
wire [1-1:0] m03_axi_arready;
wire [C_M03_AXI_ADDR_WIDTH-1:0] m03_axi_araddr;
wire [8-1:0] m03_axi_arlen;
wire [1-1:0] m03_axi_rvalid;
wire [1-1:0] m03_axi_rready;
wire [C_M03_AXI_DATA_WIDTH-1:0] m03_axi_rdata;
wire [1-1:0] m03_axi_rlast;
//AXI4 master interface m04_axi
wire [1-1:0] m04_axi_awvalid;
wire [1-1:0] m04_axi_awready;
wire [C_M04_AXI_ADDR_WIDTH-1:0] m04_axi_awaddr;
wire [8-1:0] m04_axi_awlen;
wire [1-1:0] m04_axi_wvalid;
wire [1-1:0] m04_axi_wready;
wire [C_M04_AXI_DATA_WIDTH-1:0] m04_axi_wdata;
wire [C_M04_AXI_DATA_WIDTH/8-1:0] m04_axi_wstrb;
wire [1-1:0] m04_axi_wlast;
wire [1-1:0] m04_axi_bvalid;
wire [1-1:0] m04_axi_bready;
wire [1-1:0] m04_axi_arvalid;
wire [1-1:0] m04_axi_arready;
wire [C_M04_AXI_ADDR_WIDTH-1:0] m04_axi_araddr;
wire [8-1:0] m04_axi_arlen;
wire [1-1:0] m04_axi_rvalid;
wire [1-1:0] m04_axi_rready;
wire [C_M04_AXI_DATA_WIDTH-1:0] m04_axi_rdata;
wire [1-1:0] m04_axi_rlast;
//AXI4 master interface m05_axi
wire [1-1:0] m05_axi_awvalid;
wire [1-1:0] m05_axi_awready;
wire [C_M05_AXI_ADDR_WIDTH-1:0] m05_axi_awaddr;
wire [8-1:0] m05_axi_awlen;
wire [1-1:0] m05_axi_wvalid;
wire [1-1:0] m05_axi_wready;
wire [C_M05_AXI_DATA_WIDTH-1:0] m05_axi_wdata;
wire [C_M05_AXI_DATA_WIDTH/8-1:0] m05_axi_wstrb;
wire [1-1:0] m05_axi_wlast;
wire [1-1:0] m05_axi_bvalid;
wire [1-1:0] m05_axi_bready;
wire [1-1:0] m05_axi_arvalid;
wire [1-1:0] m05_axi_arready;
wire [C_M05_AXI_ADDR_WIDTH-1:0] m05_axi_araddr;
wire [8-1:0] m05_axi_arlen;
wire [1-1:0] m05_axi_rvalid;
wire [1-1:0] m05_axi_rready;
wire [C_M05_AXI_DATA_WIDTH-1:0] m05_axi_rdata;
wire [1-1:0] m05_axi_rlast;
//AXI4 master interface m06_axi
wire [1-1:0] m06_axi_awvalid;
wire [1-1:0] m06_axi_awready;
wire [C_M06_AXI_ADDR_WIDTH-1:0] m06_axi_awaddr;
wire [8-1:0] m06_axi_awlen;
wire [1-1:0] m06_axi_wvalid;
wire [1-1:0] m06_axi_wready;
wire [C_M06_AXI_DATA_WIDTH-1:0] m06_axi_wdata;
wire [C_M06_AXI_DATA_WIDTH/8-1:0] m06_axi_wstrb;
wire [1-1:0] m06_axi_wlast;
wire [1-1:0] m06_axi_bvalid;
wire [1-1:0] m06_axi_bready;
wire [1-1:0] m06_axi_arvalid;
wire [1-1:0] m06_axi_arready;
wire [C_M06_AXI_ADDR_WIDTH-1:0] m06_axi_araddr;
wire [8-1:0] m06_axi_arlen;
wire [1-1:0] m06_axi_rvalid;
wire [1-1:0] m06_axi_rready;
wire [C_M06_AXI_DATA_WIDTH-1:0] m06_axi_rdata;
wire [1-1:0] m06_axi_rlast;
//AXI4 master interface m07_axi
wire [1-1:0] m07_axi_awvalid;
wire [1-1:0] m07_axi_awready;
wire [C_M07_AXI_ADDR_WIDTH-1:0] m07_axi_awaddr;
wire [8-1:0] m07_axi_awlen;
wire [1-1:0] m07_axi_wvalid;
wire [1-1:0] m07_axi_wready;
wire [C_M07_AXI_DATA_WIDTH-1:0] m07_axi_wdata;
wire [C_M07_AXI_DATA_WIDTH/8-1:0] m07_axi_wstrb;
wire [1-1:0] m07_axi_wlast;
wire [1-1:0] m07_axi_bvalid;
wire [1-1:0] m07_axi_bready;
wire [1-1:0] m07_axi_arvalid;
wire [1-1:0] m07_axi_arready;
wire [C_M07_AXI_ADDR_WIDTH-1:0] m07_axi_araddr;
wire [8-1:0] m07_axi_arlen;
wire [1-1:0] m07_axi_rvalid;
wire [1-1:0] m07_axi_rready;
wire [C_M07_AXI_DATA_WIDTH-1:0] m07_axi_rdata;
wire [1-1:0] m07_axi_rlast;
//AXI4 master interface m08_axi
wire [1-1:0] m08_axi_awvalid;
wire [1-1:0] m08_axi_awready;
wire [C_M08_AXI_ADDR_WIDTH-1:0] m08_axi_awaddr;
wire [8-1:0] m08_axi_awlen;
wire [1-1:0] m08_axi_wvalid;
wire [1-1:0] m08_axi_wready;
wire [C_M08_AXI_DATA_WIDTH-1:0] m08_axi_wdata;
wire [C_M08_AXI_DATA_WIDTH/8-1:0] m08_axi_wstrb;
wire [1-1:0] m08_axi_wlast;
wire [1-1:0] m08_axi_bvalid;
wire [1-1:0] m08_axi_bready;
wire [1-1:0] m08_axi_arvalid;
wire [1-1:0] m08_axi_arready;
wire [C_M08_AXI_ADDR_WIDTH-1:0] m08_axi_araddr;
wire [8-1:0] m08_axi_arlen;
wire [1-1:0] m08_axi_rvalid;
wire [1-1:0] m08_axi_rready;
wire [C_M08_AXI_DATA_WIDTH-1:0] m08_axi_rdata;
wire [1-1:0] m08_axi_rlast;
//AXI4 master interface m09_axi
wire [1-1:0] m09_axi_awvalid;
wire [1-1:0] m09_axi_awready;
wire [C_M09_AXI_ADDR_WIDTH-1:0] m09_axi_awaddr;
wire [8-1:0] m09_axi_awlen;
wire [1-1:0] m09_axi_wvalid;
wire [1-1:0] m09_axi_wready;
wire [C_M09_AXI_DATA_WIDTH-1:0] m09_axi_wdata;
wire [C_M09_AXI_DATA_WIDTH/8-1:0] m09_axi_wstrb;
wire [1-1:0] m09_axi_wlast;
wire [1-1:0] m09_axi_bvalid;
wire [1-1:0] m09_axi_bready;
wire [1-1:0] m09_axi_arvalid;
wire [1-1:0] m09_axi_arready;
wire [C_M09_AXI_ADDR_WIDTH-1:0] m09_axi_araddr;
wire [8-1:0] m09_axi_arlen;
wire [1-1:0] m09_axi_rvalid;
wire [1-1:0] m09_axi_rready;
wire [C_M09_AXI_DATA_WIDTH-1:0] m09_axi_rdata;
wire [1-1:0] m09_axi_rlast;
//AXI4 master interface m10_axi
wire [1-1:0] m10_axi_awvalid;
wire [1-1:0] m10_axi_awready;
wire [C_M10_AXI_ADDR_WIDTH-1:0] m10_axi_awaddr;
wire [8-1:0] m10_axi_awlen;
wire [1-1:0] m10_axi_wvalid;
wire [1-1:0] m10_axi_wready;
wire [C_M10_AXI_DATA_WIDTH-1:0] m10_axi_wdata;
wire [C_M10_AXI_DATA_WIDTH/8-1:0] m10_axi_wstrb;
wire [1-1:0] m10_axi_wlast;
wire [1-1:0] m10_axi_bvalid;
wire [1-1:0] m10_axi_bready;
wire [1-1:0] m10_axi_arvalid;
wire [1-1:0] m10_axi_arready;
wire [C_M10_AXI_ADDR_WIDTH-1:0] m10_axi_araddr;
wire [8-1:0] m10_axi_arlen;
wire [1-1:0] m10_axi_rvalid;
wire [1-1:0] m10_axi_rready;
wire [C_M10_AXI_DATA_WIDTH-1:0] m10_axi_rdata;
wire [1-1:0] m10_axi_rlast;
//AXI4 master interface m11_axi
wire [1-1:0] m11_axi_awvalid;
wire [1-1:0] m11_axi_awready;
wire [C_M11_AXI_ADDR_WIDTH-1:0] m11_axi_awaddr;
wire [8-1:0] m11_axi_awlen;
wire [1-1:0] m11_axi_wvalid;
wire [1-1:0] m11_axi_wready;
wire [C_M11_AXI_DATA_WIDTH-1:0] m11_axi_wdata;
wire [C_M11_AXI_DATA_WIDTH/8-1:0] m11_axi_wstrb;
wire [1-1:0] m11_axi_wlast;
wire [1-1:0] m11_axi_bvalid;
wire [1-1:0] m11_axi_bready;
wire [1-1:0] m11_axi_arvalid;
wire [1-1:0] m11_axi_arready;
wire [C_M11_AXI_ADDR_WIDTH-1:0] m11_axi_araddr;
wire [8-1:0] m11_axi_arlen;
wire [1-1:0] m11_axi_rvalid;
wire [1-1:0] m11_axi_rready;
wire [C_M11_AXI_DATA_WIDTH-1:0] m11_axi_rdata;
wire [1-1:0] m11_axi_rlast;
//AXI4 master interface m12_axi
wire [1-1:0] m12_axi_awvalid;
wire [1-1:0] m12_axi_awready;
wire [C_M12_AXI_ADDR_WIDTH-1:0] m12_axi_awaddr;
wire [8-1:0] m12_axi_awlen;
wire [1-1:0] m12_axi_wvalid;
wire [1-1:0] m12_axi_wready;
wire [C_M12_AXI_DATA_WIDTH-1:0] m12_axi_wdata;
wire [C_M12_AXI_DATA_WIDTH/8-1:0] m12_axi_wstrb;
wire [1-1:0] m12_axi_wlast;
wire [1-1:0] m12_axi_bvalid;
wire [1-1:0] m12_axi_bready;
wire [1-1:0] m12_axi_arvalid;
wire [1-1:0] m12_axi_arready;
wire [C_M12_AXI_ADDR_WIDTH-1:0] m12_axi_araddr;
wire [8-1:0] m12_axi_arlen;
wire [1-1:0] m12_axi_rvalid;
wire [1-1:0] m12_axi_rready;
wire [C_M12_AXI_DATA_WIDTH-1:0] m12_axi_rdata;
wire [1-1:0] m12_axi_rlast;
//AXI4 master interface m13_axi
wire [1-1:0] m13_axi_awvalid;
wire [1-1:0] m13_axi_awready;
wire [C_M13_AXI_ADDR_WIDTH-1:0] m13_axi_awaddr;
wire [8-1:0] m13_axi_awlen;
wire [1-1:0] m13_axi_wvalid;
wire [1-1:0] m13_axi_wready;
wire [C_M13_AXI_DATA_WIDTH-1:0] m13_axi_wdata;
wire [C_M13_AXI_DATA_WIDTH/8-1:0] m13_axi_wstrb;
wire [1-1:0] m13_axi_wlast;
wire [1-1:0] m13_axi_bvalid;
wire [1-1:0] m13_axi_bready;
wire [1-1:0] m13_axi_arvalid;
wire [1-1:0] m13_axi_arready;
wire [C_M13_AXI_ADDR_WIDTH-1:0] m13_axi_araddr;
wire [8-1:0] m13_axi_arlen;
wire [1-1:0] m13_axi_rvalid;
wire [1-1:0] m13_axi_rready;
wire [C_M13_AXI_DATA_WIDTH-1:0] m13_axi_rdata;
wire [1-1:0] m13_axi_rlast;
//AXI4 master interface m14_axi
wire [1-1:0] m14_axi_awvalid;
wire [1-1:0] m14_axi_awready;
wire [C_M14_AXI_ADDR_WIDTH-1:0] m14_axi_awaddr;
wire [8-1:0] m14_axi_awlen;
wire [1-1:0] m14_axi_wvalid;
wire [1-1:0] m14_axi_wready;
wire [C_M14_AXI_DATA_WIDTH-1:0] m14_axi_wdata;
wire [C_M14_AXI_DATA_WIDTH/8-1:0] m14_axi_wstrb;
wire [1-1:0] m14_axi_wlast;
wire [1-1:0] m14_axi_bvalid;
wire [1-1:0] m14_axi_bready;
wire [1-1:0] m14_axi_arvalid;
wire [1-1:0] m14_axi_arready;
wire [C_M14_AXI_ADDR_WIDTH-1:0] m14_axi_araddr;
wire [8-1:0] m14_axi_arlen;
wire [1-1:0] m14_axi_rvalid;
wire [1-1:0] m14_axi_rready;
wire [C_M14_AXI_DATA_WIDTH-1:0] m14_axi_rdata;
wire [1-1:0] m14_axi_rlast;
//AXI4 master interface m15_axi
wire [1-1:0] m15_axi_awvalid;
wire [1-1:0] m15_axi_awready;
wire [C_M15_AXI_ADDR_WIDTH-1:0] m15_axi_awaddr;
wire [8-1:0] m15_axi_awlen;
wire [1-1:0] m15_axi_wvalid;
wire [1-1:0] m15_axi_wready;
wire [C_M15_AXI_DATA_WIDTH-1:0] m15_axi_wdata;
wire [C_M15_AXI_DATA_WIDTH/8-1:0] m15_axi_wstrb;
wire [1-1:0] m15_axi_wlast;
wire [1-1:0] m15_axi_bvalid;
wire [1-1:0] m15_axi_bready;
wire [1-1:0] m15_axi_arvalid;
wire [1-1:0] m15_axi_arready;
wire [C_M15_AXI_ADDR_WIDTH-1:0] m15_axi_araddr;
wire [8-1:0] m15_axi_arlen;
wire [1-1:0] m15_axi_rvalid;
wire [1-1:0] m15_axi_rready;
wire [C_M15_AXI_DATA_WIDTH-1:0] m15_axi_rdata;
wire [1-1:0] m15_axi_rlast;
//AXI4 master interface m16_axi
wire [1-1:0] m16_axi_awvalid;
wire [1-1:0] m16_axi_awready;
wire [C_M16_AXI_ADDR_WIDTH-1:0] m16_axi_awaddr;
wire [8-1:0] m16_axi_awlen;
wire [1-1:0] m16_axi_wvalid;
wire [1-1:0] m16_axi_wready;
wire [C_M16_AXI_DATA_WIDTH-1:0] m16_axi_wdata;
wire [C_M16_AXI_DATA_WIDTH/8-1:0] m16_axi_wstrb;
wire [1-1:0] m16_axi_wlast;
wire [1-1:0] m16_axi_bvalid;
wire [1-1:0] m16_axi_bready;
wire [1-1:0] m16_axi_arvalid;
wire [1-1:0] m16_axi_arready;
wire [C_M16_AXI_ADDR_WIDTH-1:0] m16_axi_araddr;
wire [8-1:0] m16_axi_arlen;
wire [1-1:0] m16_axi_rvalid;
wire [1-1:0] m16_axi_rready;
wire [C_M16_AXI_DATA_WIDTH-1:0] m16_axi_rdata;
wire [1-1:0] m16_axi_rlast;
//AXI4 master interface m17_axi
wire [1-1:0] m17_axi_awvalid;
wire [1-1:0] m17_axi_awready;
wire [C_M17_AXI_ADDR_WIDTH-1:0] m17_axi_awaddr;
wire [8-1:0] m17_axi_awlen;
wire [1-1:0] m17_axi_wvalid;
wire [1-1:0] m17_axi_wready;
wire [C_M17_AXI_DATA_WIDTH-1:0] m17_axi_wdata;
wire [C_M17_AXI_DATA_WIDTH/8-1:0] m17_axi_wstrb;
wire [1-1:0] m17_axi_wlast;
wire [1-1:0] m17_axi_bvalid;
wire [1-1:0] m17_axi_bready;
wire [1-1:0] m17_axi_arvalid;
wire [1-1:0] m17_axi_arready;
wire [C_M17_AXI_ADDR_WIDTH-1:0] m17_axi_araddr;
wire [8-1:0] m17_axi_arlen;
wire [1-1:0] m17_axi_rvalid;
wire [1-1:0] m17_axi_rready;
wire [C_M17_AXI_DATA_WIDTH-1:0] m17_axi_rdata;
wire [1-1:0] m17_axi_rlast;
//AXI4 master interface m18_axi
wire [1-1:0] m18_axi_awvalid;
wire [1-1:0] m18_axi_awready;
wire [C_M18_AXI_ADDR_WIDTH-1:0] m18_axi_awaddr;
wire [8-1:0] m18_axi_awlen;
wire [1-1:0] m18_axi_wvalid;
wire [1-1:0] m18_axi_wready;
wire [C_M18_AXI_DATA_WIDTH-1:0] m18_axi_wdata;
wire [C_M18_AXI_DATA_WIDTH/8-1:0] m18_axi_wstrb;
wire [1-1:0] m18_axi_wlast;
wire [1-1:0] m18_axi_bvalid;
wire [1-1:0] m18_axi_bready;
wire [1-1:0] m18_axi_arvalid;
wire [1-1:0] m18_axi_arready;
wire [C_M18_AXI_ADDR_WIDTH-1:0] m18_axi_araddr;
wire [8-1:0] m18_axi_arlen;
wire [1-1:0] m18_axi_rvalid;
wire [1-1:0] m18_axi_rready;
wire [C_M18_AXI_DATA_WIDTH-1:0] m18_axi_rdata;
wire [1-1:0] m18_axi_rlast;
//AXI4 master interface m19_axi
wire [1-1:0] m19_axi_awvalid;
wire [1-1:0] m19_axi_awready;
wire [C_M19_AXI_ADDR_WIDTH-1:0] m19_axi_awaddr;
wire [8-1:0] m19_axi_awlen;
wire [1-1:0] m19_axi_wvalid;
wire [1-1:0] m19_axi_wready;
wire [C_M19_AXI_DATA_WIDTH-1:0] m19_axi_wdata;
wire [C_M19_AXI_DATA_WIDTH/8-1:0] m19_axi_wstrb;
wire [1-1:0] m19_axi_wlast;
wire [1-1:0] m19_axi_bvalid;
wire [1-1:0] m19_axi_bready;
wire [1-1:0] m19_axi_arvalid;
wire [1-1:0] m19_axi_arready;
wire [C_M19_AXI_ADDR_WIDTH-1:0] m19_axi_araddr;
wire [8-1:0] m19_axi_arlen;
wire [1-1:0] m19_axi_rvalid;
wire [1-1:0] m19_axi_rready;
wire [C_M19_AXI_DATA_WIDTH-1:0] m19_axi_rdata;
wire [1-1:0] m19_axi_rlast;
//AXI4 master interface m20_axi
wire [1-1:0] m20_axi_awvalid;
wire [1-1:0] m20_axi_awready;
wire [C_M20_AXI_ADDR_WIDTH-1:0] m20_axi_awaddr;
wire [8-1:0] m20_axi_awlen;
wire [1-1:0] m20_axi_wvalid;
wire [1-1:0] m20_axi_wready;
wire [C_M20_AXI_DATA_WIDTH-1:0] m20_axi_wdata;
wire [C_M20_AXI_DATA_WIDTH/8-1:0] m20_axi_wstrb;
wire [1-1:0] m20_axi_wlast;
wire [1-1:0] m20_axi_bvalid;
wire [1-1:0] m20_axi_bready;
wire [1-1:0] m20_axi_arvalid;
wire [1-1:0] m20_axi_arready;
wire [C_M20_AXI_ADDR_WIDTH-1:0] m20_axi_araddr;
wire [8-1:0] m20_axi_arlen;
wire [1-1:0] m20_axi_rvalid;
wire [1-1:0] m20_axi_rready;
wire [C_M20_AXI_DATA_WIDTH-1:0] m20_axi_rdata;
wire [1-1:0] m20_axi_rlast;
//AXI4 master interface m21_axi
wire [1-1:0] m21_axi_awvalid;
wire [1-1:0] m21_axi_awready;
wire [C_M21_AXI_ADDR_WIDTH-1:0] m21_axi_awaddr;
wire [8-1:0] m21_axi_awlen;
wire [1-1:0] m21_axi_wvalid;
wire [1-1:0] m21_axi_wready;
wire [C_M21_AXI_DATA_WIDTH-1:0] m21_axi_wdata;
wire [C_M21_AXI_DATA_WIDTH/8-1:0] m21_axi_wstrb;
wire [1-1:0] m21_axi_wlast;
wire [1-1:0] m21_axi_bvalid;
wire [1-1:0] m21_axi_bready;
wire [1-1:0] m21_axi_arvalid;
wire [1-1:0] m21_axi_arready;
wire [C_M21_AXI_ADDR_WIDTH-1:0] m21_axi_araddr;
wire [8-1:0] m21_axi_arlen;
wire [1-1:0] m21_axi_rvalid;
wire [1-1:0] m21_axi_rready;
wire [C_M21_AXI_DATA_WIDTH-1:0] m21_axi_rdata;
wire [1-1:0] m21_axi_rlast;
//AXI4 master interface m22_axi
wire [1-1:0] m22_axi_awvalid;
wire [1-1:0] m22_axi_awready;
wire [C_M22_AXI_ADDR_WIDTH-1:0] m22_axi_awaddr;
wire [8-1:0] m22_axi_awlen;
wire [1-1:0] m22_axi_wvalid;
wire [1-1:0] m22_axi_wready;
wire [C_M22_AXI_DATA_WIDTH-1:0] m22_axi_wdata;
wire [C_M22_AXI_DATA_WIDTH/8-1:0] m22_axi_wstrb;
wire [1-1:0] m22_axi_wlast;
wire [1-1:0] m22_axi_bvalid;
wire [1-1:0] m22_axi_bready;
wire [1-1:0] m22_axi_arvalid;
wire [1-1:0] m22_axi_arready;
wire [C_M22_AXI_ADDR_WIDTH-1:0] m22_axi_araddr;
wire [8-1:0] m22_axi_arlen;
wire [1-1:0] m22_axi_rvalid;
wire [1-1:0] m22_axi_rready;
wire [C_M22_AXI_DATA_WIDTH-1:0] m22_axi_rdata;
wire [1-1:0] m22_axi_rlast;
//AXI4 master interface m23_axi
wire [1-1:0] m23_axi_awvalid;
wire [1-1:0] m23_axi_awready;
wire [C_M23_AXI_ADDR_WIDTH-1:0] m23_axi_awaddr;
wire [8-1:0] m23_axi_awlen;
wire [1-1:0] m23_axi_wvalid;
wire [1-1:0] m23_axi_wready;
wire [C_M23_AXI_DATA_WIDTH-1:0] m23_axi_wdata;
wire [C_M23_AXI_DATA_WIDTH/8-1:0] m23_axi_wstrb;
wire [1-1:0] m23_axi_wlast;
wire [1-1:0] m23_axi_bvalid;
wire [1-1:0] m23_axi_bready;
wire [1-1:0] m23_axi_arvalid;
wire [1-1:0] m23_axi_arready;
wire [C_M23_AXI_ADDR_WIDTH-1:0] m23_axi_araddr;
wire [8-1:0] m23_axi_arlen;
wire [1-1:0] m23_axi_rvalid;
wire [1-1:0] m23_axi_rready;
wire [C_M23_AXI_DATA_WIDTH-1:0] m23_axi_rdata;
wire [1-1:0] m23_axi_rlast;
//AXI4 master interface m24_axi
wire [1-1:0] m24_axi_awvalid;
wire [1-1:0] m24_axi_awready;
wire [C_M24_AXI_ADDR_WIDTH-1:0] m24_axi_awaddr;
wire [8-1:0] m24_axi_awlen;
wire [1-1:0] m24_axi_wvalid;
wire [1-1:0] m24_axi_wready;
wire [C_M24_AXI_DATA_WIDTH-1:0] m24_axi_wdata;
wire [C_M24_AXI_DATA_WIDTH/8-1:0] m24_axi_wstrb;
wire [1-1:0] m24_axi_wlast;
wire [1-1:0] m24_axi_bvalid;
wire [1-1:0] m24_axi_bready;
wire [1-1:0] m24_axi_arvalid;
wire [1-1:0] m24_axi_arready;
wire [C_M24_AXI_ADDR_WIDTH-1:0] m24_axi_araddr;
wire [8-1:0] m24_axi_arlen;
wire [1-1:0] m24_axi_rvalid;
wire [1-1:0] m24_axi_rready;
wire [C_M24_AXI_DATA_WIDTH-1:0] m24_axi_rdata;
wire [1-1:0] m24_axi_rlast;
//AXI4 master interface m25_axi
wire [1-1:0] m25_axi_awvalid;
wire [1-1:0] m25_axi_awready;
wire [C_M25_AXI_ADDR_WIDTH-1:0] m25_axi_awaddr;
wire [8-1:0] m25_axi_awlen;
wire [1-1:0] m25_axi_wvalid;
wire [1-1:0] m25_axi_wready;
wire [C_M25_AXI_DATA_WIDTH-1:0] m25_axi_wdata;
wire [C_M25_AXI_DATA_WIDTH/8-1:0] m25_axi_wstrb;
wire [1-1:0] m25_axi_wlast;
wire [1-1:0] m25_axi_bvalid;
wire [1-1:0] m25_axi_bready;
wire [1-1:0] m25_axi_arvalid;
wire [1-1:0] m25_axi_arready;
wire [C_M25_AXI_ADDR_WIDTH-1:0] m25_axi_araddr;
wire [8-1:0] m25_axi_arlen;
wire [1-1:0] m25_axi_rvalid;
wire [1-1:0] m25_axi_rready;
wire [C_M25_AXI_DATA_WIDTH-1:0] m25_axi_rdata;
wire [1-1:0] m25_axi_rlast;
//AXI4 master interface m26_axi
wire [1-1:0] m26_axi_awvalid;
wire [1-1:0] m26_axi_awready;
wire [C_M26_AXI_ADDR_WIDTH-1:0] m26_axi_awaddr;
wire [8-1:0] m26_axi_awlen;
wire [1-1:0] m26_axi_wvalid;
wire [1-1:0] m26_axi_wready;
wire [C_M26_AXI_DATA_WIDTH-1:0] m26_axi_wdata;
wire [C_M26_AXI_DATA_WIDTH/8-1:0] m26_axi_wstrb;
wire [1-1:0] m26_axi_wlast;
wire [1-1:0] m26_axi_bvalid;
wire [1-1:0] m26_axi_bready;
wire [1-1:0] m26_axi_arvalid;
wire [1-1:0] m26_axi_arready;
wire [C_M26_AXI_ADDR_WIDTH-1:0] m26_axi_araddr;
wire [8-1:0] m26_axi_arlen;
wire [1-1:0] m26_axi_rvalid;
wire [1-1:0] m26_axi_rready;
wire [C_M26_AXI_DATA_WIDTH-1:0] m26_axi_rdata;
wire [1-1:0] m26_axi_rlast;
//AXI4 master interface m27_axi
wire [1-1:0] m27_axi_awvalid;
wire [1-1:0] m27_axi_awready;
wire [C_M27_AXI_ADDR_WIDTH-1:0] m27_axi_awaddr;
wire [8-1:0] m27_axi_awlen;
wire [1-1:0] m27_axi_wvalid;
wire [1-1:0] m27_axi_wready;
wire [C_M27_AXI_DATA_WIDTH-1:0] m27_axi_wdata;
wire [C_M27_AXI_DATA_WIDTH/8-1:0] m27_axi_wstrb;
wire [1-1:0] m27_axi_wlast;
wire [1-1:0] m27_axi_bvalid;
wire [1-1:0] m27_axi_bready;
wire [1-1:0] m27_axi_arvalid;
wire [1-1:0] m27_axi_arready;
wire [C_M27_AXI_ADDR_WIDTH-1:0] m27_axi_araddr;
wire [8-1:0] m27_axi_arlen;
wire [1-1:0] m27_axi_rvalid;
wire [1-1:0] m27_axi_rready;
wire [C_M27_AXI_DATA_WIDTH-1:0] m27_axi_rdata;
wire [1-1:0] m27_axi_rlast;
//AXI4 master interface m28_axi
wire [1-1:0] m28_axi_awvalid;
wire [1-1:0] m28_axi_awready;
wire [C_M28_AXI_ADDR_WIDTH-1:0] m28_axi_awaddr;
wire [8-1:0] m28_axi_awlen;
wire [1-1:0] m28_axi_wvalid;
wire [1-1:0] m28_axi_wready;
wire [C_M28_AXI_DATA_WIDTH-1:0] m28_axi_wdata;
wire [C_M28_AXI_DATA_WIDTH/8-1:0] m28_axi_wstrb;
wire [1-1:0] m28_axi_wlast;
wire [1-1:0] m28_axi_bvalid;
wire [1-1:0] m28_axi_bready;
wire [1-1:0] m28_axi_arvalid;
wire [1-1:0] m28_axi_arready;
wire [C_M28_AXI_ADDR_WIDTH-1:0] m28_axi_araddr;
wire [8-1:0] m28_axi_arlen;
wire [1-1:0] m28_axi_rvalid;
wire [1-1:0] m28_axi_rready;
wire [C_M28_AXI_DATA_WIDTH-1:0] m28_axi_rdata;
wire [1-1:0] m28_axi_rlast;
//AXI4 master interface m29_axi
wire [1-1:0] m29_axi_awvalid;
wire [1-1:0] m29_axi_awready;
wire [C_M29_AXI_ADDR_WIDTH-1:0] m29_axi_awaddr;
wire [8-1:0] m29_axi_awlen;
wire [1-1:0] m29_axi_wvalid;
wire [1-1:0] m29_axi_wready;
wire [C_M29_AXI_DATA_WIDTH-1:0] m29_axi_wdata;
wire [C_M29_AXI_DATA_WIDTH/8-1:0] m29_axi_wstrb;
wire [1-1:0] m29_axi_wlast;
wire [1-1:0] m29_axi_bvalid;
wire [1-1:0] m29_axi_bready;
wire [1-1:0] m29_axi_arvalid;
wire [1-1:0] m29_axi_arready;
wire [C_M29_AXI_ADDR_WIDTH-1:0] m29_axi_araddr;
wire [8-1:0] m29_axi_arlen;
wire [1-1:0] m29_axi_rvalid;
wire [1-1:0] m29_axi_rready;
wire [C_M29_AXI_DATA_WIDTH-1:0] m29_axi_rdata;
wire [1-1:0] m29_axi_rlast;
//AXI4 master interface m30_axi
wire [1-1:0] m30_axi_awvalid;
wire [1-1:0] m30_axi_awready;
wire [C_M30_AXI_ADDR_WIDTH-1:0] m30_axi_awaddr;
wire [8-1:0] m30_axi_awlen;
wire [1-1:0] m30_axi_wvalid;
wire [1-1:0] m30_axi_wready;
wire [C_M30_AXI_DATA_WIDTH-1:0] m30_axi_wdata;
wire [C_M30_AXI_DATA_WIDTH/8-1:0] m30_axi_wstrb;
wire [1-1:0] m30_axi_wlast;
wire [1-1:0] m30_axi_bvalid;
wire [1-1:0] m30_axi_bready;
wire [1-1:0] m30_axi_arvalid;
wire [1-1:0] m30_axi_arready;
wire [C_M30_AXI_ADDR_WIDTH-1:0] m30_axi_araddr;
wire [8-1:0] m30_axi_arlen;
wire [1-1:0] m30_axi_rvalid;
wire [1-1:0] m30_axi_rready;
wire [C_M30_AXI_DATA_WIDTH-1:0] m30_axi_rdata;
wire [1-1:0] m30_axi_rlast;
//AXI4 master interface m31_axi
wire [1-1:0] m31_axi_awvalid;
wire [1-1:0] m31_axi_awready;
wire [C_M31_AXI_ADDR_WIDTH-1:0] m31_axi_awaddr;
wire [8-1:0] m31_axi_awlen;
wire [1-1:0] m31_axi_wvalid;
wire [1-1:0] m31_axi_wready;
wire [C_M31_AXI_DATA_WIDTH-1:0] m31_axi_wdata;
wire [C_M31_AXI_DATA_WIDTH/8-1:0] m31_axi_wstrb;
wire [1-1:0] m31_axi_wlast;
wire [1-1:0] m31_axi_bvalid;
wire [1-1:0] m31_axi_bready;
wire [1-1:0] m31_axi_arvalid;
wire [1-1:0] m31_axi_arready;
wire [C_M31_AXI_ADDR_WIDTH-1:0] m31_axi_araddr;
wire [8-1:0] m31_axi_arlen;
wire [1-1:0] m31_axi_rvalid;
wire [1-1:0] m31_axi_rready;
wire [C_M31_AXI_DATA_WIDTH-1:0] m31_axi_rdata;
wire [1-1:0] m31_axi_rlast;
//AXI4LITE control signals
wire [1-1:0] s_axi_control_awvalid;
wire [1-1:0] s_axi_control_awready;
wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_awaddr;
wire [1-1:0] s_axi_control_wvalid;
wire [1-1:0] s_axi_control_wready;
wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_wdata;
wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_wstrb;
wire [1-1:0] s_axi_control_arvalid;
wire [1-1:0] s_axi_control_arready;
wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0] s_axi_control_araddr;
wire [1-1:0] s_axi_control_rvalid;
wire [1-1:0] s_axi_control_rready;
wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0] s_axi_control_rdata;
wire [2-1:0] s_axi_control_rresp;
wire [1-1:0] s_axi_control_bvalid;
wire [1-1:0] s_axi_control_bready;
wire [2-1:0] s_axi_control_bresp;
wire interrupt;

//hbm_data_file location
string file_location = "/sdb/pancg/acc/data/";

// DUT instantiation
acc_kernel #(
  .C_S_AXI_CONTROL_ADDR_WIDTH ( C_S_AXI_CONTROL_ADDR_WIDTH ),
  .C_S_AXI_CONTROL_DATA_WIDTH ( C_S_AXI_CONTROL_DATA_WIDTH ),
  .C_M00_AXI_ADDR_WIDTH       ( C_M00_AXI_ADDR_WIDTH       ),
  .C_M00_AXI_DATA_WIDTH       ( C_M00_AXI_DATA_WIDTH       ),
  .C_M01_AXI_ADDR_WIDTH       ( C_M01_AXI_ADDR_WIDTH       ),
  .C_M01_AXI_DATA_WIDTH       ( C_M01_AXI_DATA_WIDTH       ),
  .C_M02_AXI_ADDR_WIDTH       ( C_M02_AXI_ADDR_WIDTH       ),
  .C_M02_AXI_DATA_WIDTH       ( C_M02_AXI_DATA_WIDTH       ),
  .C_M03_AXI_ADDR_WIDTH       ( C_M03_AXI_ADDR_WIDTH       ),
  .C_M03_AXI_DATA_WIDTH       ( C_M03_AXI_DATA_WIDTH       ),
  .C_M04_AXI_ADDR_WIDTH       ( C_M04_AXI_ADDR_WIDTH       ),
  .C_M04_AXI_DATA_WIDTH       ( C_M04_AXI_DATA_WIDTH       ),
  .C_M05_AXI_ADDR_WIDTH       ( C_M05_AXI_ADDR_WIDTH       ),
  .C_M05_AXI_DATA_WIDTH       ( C_M05_AXI_DATA_WIDTH       ),
  .C_M06_AXI_ADDR_WIDTH       ( C_M06_AXI_ADDR_WIDTH       ),
  .C_M06_AXI_DATA_WIDTH       ( C_M06_AXI_DATA_WIDTH       ),
  .C_M07_AXI_ADDR_WIDTH       ( C_M07_AXI_ADDR_WIDTH       ),
  .C_M07_AXI_DATA_WIDTH       ( C_M07_AXI_DATA_WIDTH       ),
  .C_M08_AXI_ADDR_WIDTH       ( C_M08_AXI_ADDR_WIDTH       ),
  .C_M08_AXI_DATA_WIDTH       ( C_M08_AXI_DATA_WIDTH       ),
  .C_M09_AXI_ADDR_WIDTH       ( C_M09_AXI_ADDR_WIDTH       ),
  .C_M09_AXI_DATA_WIDTH       ( C_M09_AXI_DATA_WIDTH       ),
  .C_M10_AXI_ADDR_WIDTH       ( C_M10_AXI_ADDR_WIDTH       ),
  .C_M10_AXI_DATA_WIDTH       ( C_M10_AXI_DATA_WIDTH       ),
  .C_M11_AXI_ADDR_WIDTH       ( C_M11_AXI_ADDR_WIDTH       ),
  .C_M11_AXI_DATA_WIDTH       ( C_M11_AXI_DATA_WIDTH       ),
  .C_M12_AXI_ADDR_WIDTH       ( C_M12_AXI_ADDR_WIDTH       ),
  .C_M12_AXI_DATA_WIDTH       ( C_M12_AXI_DATA_WIDTH       ),
  .C_M13_AXI_ADDR_WIDTH       ( C_M13_AXI_ADDR_WIDTH       ),
  .C_M13_AXI_DATA_WIDTH       ( C_M13_AXI_DATA_WIDTH       ),
  .C_M14_AXI_ADDR_WIDTH       ( C_M14_AXI_ADDR_WIDTH       ),
  .C_M14_AXI_DATA_WIDTH       ( C_M14_AXI_DATA_WIDTH       ),
  .C_M15_AXI_ADDR_WIDTH       ( C_M15_AXI_ADDR_WIDTH       ),
  .C_M15_AXI_DATA_WIDTH       ( C_M15_AXI_DATA_WIDTH       ),
  .C_M16_AXI_ADDR_WIDTH       ( C_M16_AXI_ADDR_WIDTH       ),
  .C_M16_AXI_DATA_WIDTH       ( C_M16_AXI_DATA_WIDTH       ),
  .C_M17_AXI_ADDR_WIDTH       ( C_M17_AXI_ADDR_WIDTH       ),
  .C_M17_AXI_DATA_WIDTH       ( C_M17_AXI_DATA_WIDTH       ),
  .C_M18_AXI_ADDR_WIDTH       ( C_M18_AXI_ADDR_WIDTH       ),
  .C_M18_AXI_DATA_WIDTH       ( C_M18_AXI_DATA_WIDTH       ),
  .C_M19_AXI_ADDR_WIDTH       ( C_M19_AXI_ADDR_WIDTH       ),
  .C_M19_AXI_DATA_WIDTH       ( C_M19_AXI_DATA_WIDTH       ),
  .C_M20_AXI_ADDR_WIDTH       ( C_M20_AXI_ADDR_WIDTH       ),
  .C_M20_AXI_DATA_WIDTH       ( C_M20_AXI_DATA_WIDTH       ),
  .C_M21_AXI_ADDR_WIDTH       ( C_M21_AXI_ADDR_WIDTH       ),
  .C_M21_AXI_DATA_WIDTH       ( C_M21_AXI_DATA_WIDTH       ),
  .C_M22_AXI_ADDR_WIDTH       ( C_M22_AXI_ADDR_WIDTH       ),
  .C_M22_AXI_DATA_WIDTH       ( C_M22_AXI_DATA_WIDTH       ),
  .C_M23_AXI_ADDR_WIDTH       ( C_M23_AXI_ADDR_WIDTH       ),
  .C_M23_AXI_DATA_WIDTH       ( C_M23_AXI_DATA_WIDTH       ),
  .C_M24_AXI_ADDR_WIDTH       ( C_M24_AXI_ADDR_WIDTH       ),
  .C_M24_AXI_DATA_WIDTH       ( C_M24_AXI_DATA_WIDTH       ),
  .C_M25_AXI_ADDR_WIDTH       ( C_M25_AXI_ADDR_WIDTH       ),
  .C_M25_AXI_DATA_WIDTH       ( C_M25_AXI_DATA_WIDTH       ),
  .C_M26_AXI_ADDR_WIDTH       ( C_M26_AXI_ADDR_WIDTH       ),
  .C_M26_AXI_DATA_WIDTH       ( C_M26_AXI_DATA_WIDTH       ),
  .C_M27_AXI_ADDR_WIDTH       ( C_M27_AXI_ADDR_WIDTH       ),
  .C_M27_AXI_DATA_WIDTH       ( C_M27_AXI_DATA_WIDTH       ),
  .C_M28_AXI_ADDR_WIDTH       ( C_M28_AXI_ADDR_WIDTH       ),
  .C_M28_AXI_DATA_WIDTH       ( C_M28_AXI_DATA_WIDTH       ),
  .C_M29_AXI_ADDR_WIDTH       ( C_M29_AXI_ADDR_WIDTH       ),
  .C_M29_AXI_DATA_WIDTH       ( C_M29_AXI_DATA_WIDTH       ),
  .C_M30_AXI_ADDR_WIDTH       ( C_M30_AXI_ADDR_WIDTH       ),
  .C_M30_AXI_DATA_WIDTH       ( C_M30_AXI_DATA_WIDTH       ),
  .C_M31_AXI_ADDR_WIDTH       ( C_M31_AXI_ADDR_WIDTH       ),
  .C_M31_AXI_DATA_WIDTH       ( C_M31_AXI_DATA_WIDTH       )
)
inst_dut (
  .ap_clk                ( ap_clk                ),
  .ap_rst_n              ( ap_rst_n              ),
  .m00_axi_awvalid       ( m00_axi_awvalid       ),
  .m00_axi_awready       ( m00_axi_awready       ),
  .m00_axi_awaddr        ( m00_axi_awaddr        ),
  .m00_axi_awlen         ( m00_axi_awlen         ),
  .m00_axi_wvalid        ( m00_axi_wvalid        ),
  .m00_axi_wready        ( m00_axi_wready        ),
  .m00_axi_wdata         ( m00_axi_wdata         ),
  .m00_axi_wstrb         ( m00_axi_wstrb         ),
  .m00_axi_wlast         ( m00_axi_wlast         ),
  .m00_axi_bvalid        ( m00_axi_bvalid        ),
  .m00_axi_bready        ( m00_axi_bready        ),
  .m00_axi_arvalid       ( m00_axi_arvalid       ),
  .m00_axi_arready       ( m00_axi_arready       ),
  .m00_axi_araddr        ( m00_axi_araddr        ),
  .m00_axi_arlen         ( m00_axi_arlen         ),
  .m00_axi_rvalid        ( m00_axi_rvalid        ),
  .m00_axi_rready        ( m00_axi_rready        ),
  .m00_axi_rdata         ( m00_axi_rdata         ),
  .m00_axi_rlast         ( m00_axi_rlast         ),
  .m01_axi_awvalid       ( m01_axi_awvalid       ),
  .m01_axi_awready       ( m01_axi_awready       ),
  .m01_axi_awaddr        ( m01_axi_awaddr        ),
  .m01_axi_awlen         ( m01_axi_awlen         ),
  .m01_axi_wvalid        ( m01_axi_wvalid        ),
  .m01_axi_wready        ( m01_axi_wready        ),
  .m01_axi_wdata         ( m01_axi_wdata         ),
  .m01_axi_wstrb         ( m01_axi_wstrb         ),
  .m01_axi_wlast         ( m01_axi_wlast         ),
  .m01_axi_bvalid        ( m01_axi_bvalid        ),
  .m01_axi_bready        ( m01_axi_bready        ),
  .m01_axi_arvalid       ( m01_axi_arvalid       ),
  .m01_axi_arready       ( m01_axi_arready       ),
  .m01_axi_araddr        ( m01_axi_araddr        ),
  .m01_axi_arlen         ( m01_axi_arlen         ),
  .m01_axi_rvalid        ( m01_axi_rvalid        ),
  .m01_axi_rready        ( m01_axi_rready        ),
  .m01_axi_rdata         ( m01_axi_rdata         ),
  .m01_axi_rlast         ( m01_axi_rlast         ),
  .m02_axi_awvalid       ( m02_axi_awvalid       ),
  .m02_axi_awready       ( m02_axi_awready       ),
  .m02_axi_awaddr        ( m02_axi_awaddr        ),
  .m02_axi_awlen         ( m02_axi_awlen         ),
  .m02_axi_wvalid        ( m02_axi_wvalid        ),
  .m02_axi_wready        ( m02_axi_wready        ),
  .m02_axi_wdata         ( m02_axi_wdata         ),
  .m02_axi_wstrb         ( m02_axi_wstrb         ),
  .m02_axi_wlast         ( m02_axi_wlast         ),
  .m02_axi_bvalid        ( m02_axi_bvalid        ),
  .m02_axi_bready        ( m02_axi_bready        ),
  .m02_axi_arvalid       ( m02_axi_arvalid       ),
  .m02_axi_arready       ( m02_axi_arready       ),
  .m02_axi_araddr        ( m02_axi_araddr        ),
  .m02_axi_arlen         ( m02_axi_arlen         ),
  .m02_axi_rvalid        ( m02_axi_rvalid        ),
  .m02_axi_rready        ( m02_axi_rready        ),
  .m02_axi_rdata         ( m02_axi_rdata         ),
  .m02_axi_rlast         ( m02_axi_rlast         ),
  .m03_axi_awvalid       ( m03_axi_awvalid       ),
  .m03_axi_awready       ( m03_axi_awready       ),
  .m03_axi_awaddr        ( m03_axi_awaddr        ),
  .m03_axi_awlen         ( m03_axi_awlen         ),
  .m03_axi_wvalid        ( m03_axi_wvalid        ),
  .m03_axi_wready        ( m03_axi_wready        ),
  .m03_axi_wdata         ( m03_axi_wdata         ),
  .m03_axi_wstrb         ( m03_axi_wstrb         ),
  .m03_axi_wlast         ( m03_axi_wlast         ),
  .m03_axi_bvalid        ( m03_axi_bvalid        ),
  .m03_axi_bready        ( m03_axi_bready        ),
  .m03_axi_arvalid       ( m03_axi_arvalid       ),
  .m03_axi_arready       ( m03_axi_arready       ),
  .m03_axi_araddr        ( m03_axi_araddr        ),
  .m03_axi_arlen         ( m03_axi_arlen         ),
  .m03_axi_rvalid        ( m03_axi_rvalid        ),
  .m03_axi_rready        ( m03_axi_rready        ),
  .m03_axi_rdata         ( m03_axi_rdata         ),
  .m03_axi_rlast         ( m03_axi_rlast         ),
  .m04_axi_awvalid       ( m04_axi_awvalid       ),
  .m04_axi_awready       ( m04_axi_awready       ),
  .m04_axi_awaddr        ( m04_axi_awaddr        ),
  .m04_axi_awlen         ( m04_axi_awlen         ),
  .m04_axi_wvalid        ( m04_axi_wvalid        ),
  .m04_axi_wready        ( m04_axi_wready        ),
  .m04_axi_wdata         ( m04_axi_wdata         ),
  .m04_axi_wstrb         ( m04_axi_wstrb         ),
  .m04_axi_wlast         ( m04_axi_wlast         ),
  .m04_axi_bvalid        ( m04_axi_bvalid        ),
  .m04_axi_bready        ( m04_axi_bready        ),
  .m04_axi_arvalid       ( m04_axi_arvalid       ),
  .m04_axi_arready       ( m04_axi_arready       ),
  .m04_axi_araddr        ( m04_axi_araddr        ),
  .m04_axi_arlen         ( m04_axi_arlen         ),
  .m04_axi_rvalid        ( m04_axi_rvalid        ),
  .m04_axi_rready        ( m04_axi_rready        ),
  .m04_axi_rdata         ( m04_axi_rdata         ),
  .m04_axi_rlast         ( m04_axi_rlast         ),
  .m05_axi_awvalid       ( m05_axi_awvalid       ),
  .m05_axi_awready       ( m05_axi_awready       ),
  .m05_axi_awaddr        ( m05_axi_awaddr        ),
  .m05_axi_awlen         ( m05_axi_awlen         ),
  .m05_axi_wvalid        ( m05_axi_wvalid        ),
  .m05_axi_wready        ( m05_axi_wready        ),
  .m05_axi_wdata         ( m05_axi_wdata         ),
  .m05_axi_wstrb         ( m05_axi_wstrb         ),
  .m05_axi_wlast         ( m05_axi_wlast         ),
  .m05_axi_bvalid        ( m05_axi_bvalid        ),
  .m05_axi_bready        ( m05_axi_bready        ),
  .m05_axi_arvalid       ( m05_axi_arvalid       ),
  .m05_axi_arready       ( m05_axi_arready       ),
  .m05_axi_araddr        ( m05_axi_araddr        ),
  .m05_axi_arlen         ( m05_axi_arlen         ),
  .m05_axi_rvalid        ( m05_axi_rvalid        ),
  .m05_axi_rready        ( m05_axi_rready        ),
  .m05_axi_rdata         ( m05_axi_rdata         ),
  .m05_axi_rlast         ( m05_axi_rlast         ),
  .m06_axi_awvalid       ( m06_axi_awvalid       ),
  .m06_axi_awready       ( m06_axi_awready       ),
  .m06_axi_awaddr        ( m06_axi_awaddr        ),
  .m06_axi_awlen         ( m06_axi_awlen         ),
  .m06_axi_wvalid        ( m06_axi_wvalid        ),
  .m06_axi_wready        ( m06_axi_wready        ),
  .m06_axi_wdata         ( m06_axi_wdata         ),
  .m06_axi_wstrb         ( m06_axi_wstrb         ),
  .m06_axi_wlast         ( m06_axi_wlast         ),
  .m06_axi_bvalid        ( m06_axi_bvalid        ),
  .m06_axi_bready        ( m06_axi_bready        ),
  .m06_axi_arvalid       ( m06_axi_arvalid       ),
  .m06_axi_arready       ( m06_axi_arready       ),
  .m06_axi_araddr        ( m06_axi_araddr        ),
  .m06_axi_arlen         ( m06_axi_arlen         ),
  .m06_axi_rvalid        ( m06_axi_rvalid        ),
  .m06_axi_rready        ( m06_axi_rready        ),
  .m06_axi_rdata         ( m06_axi_rdata         ),
  .m06_axi_rlast         ( m06_axi_rlast         ),
  .m07_axi_awvalid       ( m07_axi_awvalid       ),
  .m07_axi_awready       ( m07_axi_awready       ),
  .m07_axi_awaddr        ( m07_axi_awaddr        ),
  .m07_axi_awlen         ( m07_axi_awlen         ),
  .m07_axi_wvalid        ( m07_axi_wvalid        ),
  .m07_axi_wready        ( m07_axi_wready        ),
  .m07_axi_wdata         ( m07_axi_wdata         ),
  .m07_axi_wstrb         ( m07_axi_wstrb         ),
  .m07_axi_wlast         ( m07_axi_wlast         ),
  .m07_axi_bvalid        ( m07_axi_bvalid        ),
  .m07_axi_bready        ( m07_axi_bready        ),
  .m07_axi_arvalid       ( m07_axi_arvalid       ),
  .m07_axi_arready       ( m07_axi_arready       ),
  .m07_axi_araddr        ( m07_axi_araddr        ),
  .m07_axi_arlen         ( m07_axi_arlen         ),
  .m07_axi_rvalid        ( m07_axi_rvalid        ),
  .m07_axi_rready        ( m07_axi_rready        ),
  .m07_axi_rdata         ( m07_axi_rdata         ),
  .m07_axi_rlast         ( m07_axi_rlast         ),
  .m08_axi_awvalid       ( m08_axi_awvalid       ),
  .m08_axi_awready       ( m08_axi_awready       ),
  .m08_axi_awaddr        ( m08_axi_awaddr        ),
  .m08_axi_awlen         ( m08_axi_awlen         ),
  .m08_axi_wvalid        ( m08_axi_wvalid        ),
  .m08_axi_wready        ( m08_axi_wready        ),
  .m08_axi_wdata         ( m08_axi_wdata         ),
  .m08_axi_wstrb         ( m08_axi_wstrb         ),
  .m08_axi_wlast         ( m08_axi_wlast         ),
  .m08_axi_bvalid        ( m08_axi_bvalid        ),
  .m08_axi_bready        ( m08_axi_bready        ),
  .m08_axi_arvalid       ( m08_axi_arvalid       ),
  .m08_axi_arready       ( m08_axi_arready       ),
  .m08_axi_araddr        ( m08_axi_araddr        ),
  .m08_axi_arlen         ( m08_axi_arlen         ),
  .m08_axi_rvalid        ( m08_axi_rvalid        ),
  .m08_axi_rready        ( m08_axi_rready        ),
  .m08_axi_rdata         ( m08_axi_rdata         ),
  .m08_axi_rlast         ( m08_axi_rlast         ),
  .m09_axi_awvalid       ( m09_axi_awvalid       ),
  .m09_axi_awready       ( m09_axi_awready       ),
  .m09_axi_awaddr        ( m09_axi_awaddr        ),
  .m09_axi_awlen         ( m09_axi_awlen         ),
  .m09_axi_wvalid        ( m09_axi_wvalid        ),
  .m09_axi_wready        ( m09_axi_wready        ),
  .m09_axi_wdata         ( m09_axi_wdata         ),
  .m09_axi_wstrb         ( m09_axi_wstrb         ),
  .m09_axi_wlast         ( m09_axi_wlast         ),
  .m09_axi_bvalid        ( m09_axi_bvalid        ),
  .m09_axi_bready        ( m09_axi_bready        ),
  .m09_axi_arvalid       ( m09_axi_arvalid       ),
  .m09_axi_arready       ( m09_axi_arready       ),
  .m09_axi_araddr        ( m09_axi_araddr        ),
  .m09_axi_arlen         ( m09_axi_arlen         ),
  .m09_axi_rvalid        ( m09_axi_rvalid        ),
  .m09_axi_rready        ( m09_axi_rready        ),
  .m09_axi_rdata         ( m09_axi_rdata         ),
  .m09_axi_rlast         ( m09_axi_rlast         ),
  .m10_axi_awvalid       ( m10_axi_awvalid       ),
  .m10_axi_awready       ( m10_axi_awready       ),
  .m10_axi_awaddr        ( m10_axi_awaddr        ),
  .m10_axi_awlen         ( m10_axi_awlen         ),
  .m10_axi_wvalid        ( m10_axi_wvalid        ),
  .m10_axi_wready        ( m10_axi_wready        ),
  .m10_axi_wdata         ( m10_axi_wdata         ),
  .m10_axi_wstrb         ( m10_axi_wstrb         ),
  .m10_axi_wlast         ( m10_axi_wlast         ),
  .m10_axi_bvalid        ( m10_axi_bvalid        ),
  .m10_axi_bready        ( m10_axi_bready        ),
  .m10_axi_arvalid       ( m10_axi_arvalid       ),
  .m10_axi_arready       ( m10_axi_arready       ),
  .m10_axi_araddr        ( m10_axi_araddr        ),
  .m10_axi_arlen         ( m10_axi_arlen         ),
  .m10_axi_rvalid        ( m10_axi_rvalid        ),
  .m10_axi_rready        ( m10_axi_rready        ),
  .m10_axi_rdata         ( m10_axi_rdata         ),
  .m10_axi_rlast         ( m10_axi_rlast         ),
  .m11_axi_awvalid       ( m11_axi_awvalid       ),
  .m11_axi_awready       ( m11_axi_awready       ),
  .m11_axi_awaddr        ( m11_axi_awaddr        ),
  .m11_axi_awlen         ( m11_axi_awlen         ),
  .m11_axi_wvalid        ( m11_axi_wvalid        ),
  .m11_axi_wready        ( m11_axi_wready        ),
  .m11_axi_wdata         ( m11_axi_wdata         ),
  .m11_axi_wstrb         ( m11_axi_wstrb         ),
  .m11_axi_wlast         ( m11_axi_wlast         ),
  .m11_axi_bvalid        ( m11_axi_bvalid        ),
  .m11_axi_bready        ( m11_axi_bready        ),
  .m11_axi_arvalid       ( m11_axi_arvalid       ),
  .m11_axi_arready       ( m11_axi_arready       ),
  .m11_axi_araddr        ( m11_axi_araddr        ),
  .m11_axi_arlen         ( m11_axi_arlen         ),
  .m11_axi_rvalid        ( m11_axi_rvalid        ),
  .m11_axi_rready        ( m11_axi_rready        ),
  .m11_axi_rdata         ( m11_axi_rdata         ),
  .m11_axi_rlast         ( m11_axi_rlast         ),
  .m12_axi_awvalid       ( m12_axi_awvalid       ),
  .m12_axi_awready       ( m12_axi_awready       ),
  .m12_axi_awaddr        ( m12_axi_awaddr        ),
  .m12_axi_awlen         ( m12_axi_awlen         ),
  .m12_axi_wvalid        ( m12_axi_wvalid        ),
  .m12_axi_wready        ( m12_axi_wready        ),
  .m12_axi_wdata         ( m12_axi_wdata         ),
  .m12_axi_wstrb         ( m12_axi_wstrb         ),
  .m12_axi_wlast         ( m12_axi_wlast         ),
  .m12_axi_bvalid        ( m12_axi_bvalid        ),
  .m12_axi_bready        ( m12_axi_bready        ),
  .m12_axi_arvalid       ( m12_axi_arvalid       ),
  .m12_axi_arready       ( m12_axi_arready       ),
  .m12_axi_araddr        ( m12_axi_araddr        ),
  .m12_axi_arlen         ( m12_axi_arlen         ),
  .m12_axi_rvalid        ( m12_axi_rvalid        ),
  .m12_axi_rready        ( m12_axi_rready        ),
  .m12_axi_rdata         ( m12_axi_rdata         ),
  .m12_axi_rlast         ( m12_axi_rlast         ),
  .m13_axi_awvalid       ( m13_axi_awvalid       ),
  .m13_axi_awready       ( m13_axi_awready       ),
  .m13_axi_awaddr        ( m13_axi_awaddr        ),
  .m13_axi_awlen         ( m13_axi_awlen         ),
  .m13_axi_wvalid        ( m13_axi_wvalid        ),
  .m13_axi_wready        ( m13_axi_wready        ),
  .m13_axi_wdata         ( m13_axi_wdata         ),
  .m13_axi_wstrb         ( m13_axi_wstrb         ),
  .m13_axi_wlast         ( m13_axi_wlast         ),
  .m13_axi_bvalid        ( m13_axi_bvalid        ),
  .m13_axi_bready        ( m13_axi_bready        ),
  .m13_axi_arvalid       ( m13_axi_arvalid       ),
  .m13_axi_arready       ( m13_axi_arready       ),
  .m13_axi_araddr        ( m13_axi_araddr        ),
  .m13_axi_arlen         ( m13_axi_arlen         ),
  .m13_axi_rvalid        ( m13_axi_rvalid        ),
  .m13_axi_rready        ( m13_axi_rready        ),
  .m13_axi_rdata         ( m13_axi_rdata         ),
  .m13_axi_rlast         ( m13_axi_rlast         ),
  .m14_axi_awvalid       ( m14_axi_awvalid       ),
  .m14_axi_awready       ( m14_axi_awready       ),
  .m14_axi_awaddr        ( m14_axi_awaddr        ),
  .m14_axi_awlen         ( m14_axi_awlen         ),
  .m14_axi_wvalid        ( m14_axi_wvalid        ),
  .m14_axi_wready        ( m14_axi_wready        ),
  .m14_axi_wdata         ( m14_axi_wdata         ),
  .m14_axi_wstrb         ( m14_axi_wstrb         ),
  .m14_axi_wlast         ( m14_axi_wlast         ),
  .m14_axi_bvalid        ( m14_axi_bvalid        ),
  .m14_axi_bready        ( m14_axi_bready        ),
  .m14_axi_arvalid       ( m14_axi_arvalid       ),
  .m14_axi_arready       ( m14_axi_arready       ),
  .m14_axi_araddr        ( m14_axi_araddr        ),
  .m14_axi_arlen         ( m14_axi_arlen         ),
  .m14_axi_rvalid        ( m14_axi_rvalid        ),
  .m14_axi_rready        ( m14_axi_rready        ),
  .m14_axi_rdata         ( m14_axi_rdata         ),
  .m14_axi_rlast         ( m14_axi_rlast         ),
  .m15_axi_awvalid       ( m15_axi_awvalid       ),
  .m15_axi_awready       ( m15_axi_awready       ),
  .m15_axi_awaddr        ( m15_axi_awaddr        ),
  .m15_axi_awlen         ( m15_axi_awlen         ),
  .m15_axi_wvalid        ( m15_axi_wvalid        ),
  .m15_axi_wready        ( m15_axi_wready        ),
  .m15_axi_wdata         ( m15_axi_wdata         ),
  .m15_axi_wstrb         ( m15_axi_wstrb         ),
  .m15_axi_wlast         ( m15_axi_wlast         ),
  .m15_axi_bvalid        ( m15_axi_bvalid        ),
  .m15_axi_bready        ( m15_axi_bready        ),
  .m15_axi_arvalid       ( m15_axi_arvalid       ),
  .m15_axi_arready       ( m15_axi_arready       ),
  .m15_axi_araddr        ( m15_axi_araddr        ),
  .m15_axi_arlen         ( m15_axi_arlen         ),
  .m15_axi_rvalid        ( m15_axi_rvalid        ),
  .m15_axi_rready        ( m15_axi_rready        ),
  .m15_axi_rdata         ( m15_axi_rdata         ),
  .m15_axi_rlast         ( m15_axi_rlast         ),
  .m16_axi_awvalid       ( m16_axi_awvalid       ),
  .m16_axi_awready       ( m16_axi_awready       ),
  .m16_axi_awaddr        ( m16_axi_awaddr        ),
  .m16_axi_awlen         ( m16_axi_awlen         ),
  .m16_axi_wvalid        ( m16_axi_wvalid        ),
  .m16_axi_wready        ( m16_axi_wready        ),
  .m16_axi_wdata         ( m16_axi_wdata         ),
  .m16_axi_wstrb         ( m16_axi_wstrb         ),
  .m16_axi_wlast         ( m16_axi_wlast         ),
  .m16_axi_bvalid        ( m16_axi_bvalid        ),
  .m16_axi_bready        ( m16_axi_bready        ),
  .m16_axi_arvalid       ( m16_axi_arvalid       ),
  .m16_axi_arready       ( m16_axi_arready       ),
  .m16_axi_araddr        ( m16_axi_araddr        ),
  .m16_axi_arlen         ( m16_axi_arlen         ),
  .m16_axi_rvalid        ( m16_axi_rvalid        ),
  .m16_axi_rready        ( m16_axi_rready        ),
  .m16_axi_rdata         ( m16_axi_rdata         ),
  .m16_axi_rlast         ( m16_axi_rlast         ),
  .m17_axi_awvalid       ( m17_axi_awvalid       ),
  .m17_axi_awready       ( m17_axi_awready       ),
  .m17_axi_awaddr        ( m17_axi_awaddr        ),
  .m17_axi_awlen         ( m17_axi_awlen         ),
  .m17_axi_wvalid        ( m17_axi_wvalid        ),
  .m17_axi_wready        ( m17_axi_wready        ),
  .m17_axi_wdata         ( m17_axi_wdata         ),
  .m17_axi_wstrb         ( m17_axi_wstrb         ),
  .m17_axi_wlast         ( m17_axi_wlast         ),
  .m17_axi_bvalid        ( m17_axi_bvalid        ),
  .m17_axi_bready        ( m17_axi_bready        ),
  .m17_axi_arvalid       ( m17_axi_arvalid       ),
  .m17_axi_arready       ( m17_axi_arready       ),
  .m17_axi_araddr        ( m17_axi_araddr        ),
  .m17_axi_arlen         ( m17_axi_arlen         ),
  .m17_axi_rvalid        ( m17_axi_rvalid        ),
  .m17_axi_rready        ( m17_axi_rready        ),
  .m17_axi_rdata         ( m17_axi_rdata         ),
  .m17_axi_rlast         ( m17_axi_rlast         ),
  .m18_axi_awvalid       ( m18_axi_awvalid       ),
  .m18_axi_awready       ( m18_axi_awready       ),
  .m18_axi_awaddr        ( m18_axi_awaddr        ),
  .m18_axi_awlen         ( m18_axi_awlen         ),
  .m18_axi_wvalid        ( m18_axi_wvalid        ),
  .m18_axi_wready        ( m18_axi_wready        ),
  .m18_axi_wdata         ( m18_axi_wdata         ),
  .m18_axi_wstrb         ( m18_axi_wstrb         ),
  .m18_axi_wlast         ( m18_axi_wlast         ),
  .m18_axi_bvalid        ( m18_axi_bvalid        ),
  .m18_axi_bready        ( m18_axi_bready        ),
  .m18_axi_arvalid       ( m18_axi_arvalid       ),
  .m18_axi_arready       ( m18_axi_arready       ),
  .m18_axi_araddr        ( m18_axi_araddr        ),
  .m18_axi_arlen         ( m18_axi_arlen         ),
  .m18_axi_rvalid        ( m18_axi_rvalid        ),
  .m18_axi_rready        ( m18_axi_rready        ),
  .m18_axi_rdata         ( m18_axi_rdata         ),
  .m18_axi_rlast         ( m18_axi_rlast         ),
  .m19_axi_awvalid       ( m19_axi_awvalid       ),
  .m19_axi_awready       ( m19_axi_awready       ),
  .m19_axi_awaddr        ( m19_axi_awaddr        ),
  .m19_axi_awlen         ( m19_axi_awlen         ),
  .m19_axi_wvalid        ( m19_axi_wvalid        ),
  .m19_axi_wready        ( m19_axi_wready        ),
  .m19_axi_wdata         ( m19_axi_wdata         ),
  .m19_axi_wstrb         ( m19_axi_wstrb         ),
  .m19_axi_wlast         ( m19_axi_wlast         ),
  .m19_axi_bvalid        ( m19_axi_bvalid        ),
  .m19_axi_bready        ( m19_axi_bready        ),
  .m19_axi_arvalid       ( m19_axi_arvalid       ),
  .m19_axi_arready       ( m19_axi_arready       ),
  .m19_axi_araddr        ( m19_axi_araddr        ),
  .m19_axi_arlen         ( m19_axi_arlen         ),
  .m19_axi_rvalid        ( m19_axi_rvalid        ),
  .m19_axi_rready        ( m19_axi_rready        ),
  .m19_axi_rdata         ( m19_axi_rdata         ),
  .m19_axi_rlast         ( m19_axi_rlast         ),
  .m20_axi_awvalid       ( m20_axi_awvalid       ),
  .m20_axi_awready       ( m20_axi_awready       ),
  .m20_axi_awaddr        ( m20_axi_awaddr        ),
  .m20_axi_awlen         ( m20_axi_awlen         ),
  .m20_axi_wvalid        ( m20_axi_wvalid        ),
  .m20_axi_wready        ( m20_axi_wready        ),
  .m20_axi_wdata         ( m20_axi_wdata         ),
  .m20_axi_wstrb         ( m20_axi_wstrb         ),
  .m20_axi_wlast         ( m20_axi_wlast         ),
  .m20_axi_bvalid        ( m20_axi_bvalid        ),
  .m20_axi_bready        ( m20_axi_bready        ),
  .m20_axi_arvalid       ( m20_axi_arvalid       ),
  .m20_axi_arready       ( m20_axi_arready       ),
  .m20_axi_araddr        ( m20_axi_araddr        ),
  .m20_axi_arlen         ( m20_axi_arlen         ),
  .m20_axi_rvalid        ( m20_axi_rvalid        ),
  .m20_axi_rready        ( m20_axi_rready        ),
  .m20_axi_rdata         ( m20_axi_rdata         ),
  .m20_axi_rlast         ( m20_axi_rlast         ),
  .m21_axi_awvalid       ( m21_axi_awvalid       ),
  .m21_axi_awready       ( m21_axi_awready       ),
  .m21_axi_awaddr        ( m21_axi_awaddr        ),
  .m21_axi_awlen         ( m21_axi_awlen         ),
  .m21_axi_wvalid        ( m21_axi_wvalid        ),
  .m21_axi_wready        ( m21_axi_wready        ),
  .m21_axi_wdata         ( m21_axi_wdata         ),
  .m21_axi_wstrb         ( m21_axi_wstrb         ),
  .m21_axi_wlast         ( m21_axi_wlast         ),
  .m21_axi_bvalid        ( m21_axi_bvalid        ),
  .m21_axi_bready        ( m21_axi_bready        ),
  .m21_axi_arvalid       ( m21_axi_arvalid       ),
  .m21_axi_arready       ( m21_axi_arready       ),
  .m21_axi_araddr        ( m21_axi_araddr        ),
  .m21_axi_arlen         ( m21_axi_arlen         ),
  .m21_axi_rvalid        ( m21_axi_rvalid        ),
  .m21_axi_rready        ( m21_axi_rready        ),
  .m21_axi_rdata         ( m21_axi_rdata         ),
  .m21_axi_rlast         ( m21_axi_rlast         ),
  .m22_axi_awvalid       ( m22_axi_awvalid       ),
  .m22_axi_awready       ( m22_axi_awready       ),
  .m22_axi_awaddr        ( m22_axi_awaddr        ),
  .m22_axi_awlen         ( m22_axi_awlen         ),
  .m22_axi_wvalid        ( m22_axi_wvalid        ),
  .m22_axi_wready        ( m22_axi_wready        ),
  .m22_axi_wdata         ( m22_axi_wdata         ),
  .m22_axi_wstrb         ( m22_axi_wstrb         ),
  .m22_axi_wlast         ( m22_axi_wlast         ),
  .m22_axi_bvalid        ( m22_axi_bvalid        ),
  .m22_axi_bready        ( m22_axi_bready        ),
  .m22_axi_arvalid       ( m22_axi_arvalid       ),
  .m22_axi_arready       ( m22_axi_arready       ),
  .m22_axi_araddr        ( m22_axi_araddr        ),
  .m22_axi_arlen         ( m22_axi_arlen         ),
  .m22_axi_rvalid        ( m22_axi_rvalid        ),
  .m22_axi_rready        ( m22_axi_rready        ),
  .m22_axi_rdata         ( m22_axi_rdata         ),
  .m22_axi_rlast         ( m22_axi_rlast         ),
  .m23_axi_awvalid       ( m23_axi_awvalid       ),
  .m23_axi_awready       ( m23_axi_awready       ),
  .m23_axi_awaddr        ( m23_axi_awaddr        ),
  .m23_axi_awlen         ( m23_axi_awlen         ),
  .m23_axi_wvalid        ( m23_axi_wvalid        ),
  .m23_axi_wready        ( m23_axi_wready        ),
  .m23_axi_wdata         ( m23_axi_wdata         ),
  .m23_axi_wstrb         ( m23_axi_wstrb         ),
  .m23_axi_wlast         ( m23_axi_wlast         ),
  .m23_axi_bvalid        ( m23_axi_bvalid        ),
  .m23_axi_bready        ( m23_axi_bready        ),
  .m23_axi_arvalid       ( m23_axi_arvalid       ),
  .m23_axi_arready       ( m23_axi_arready       ),
  .m23_axi_araddr        ( m23_axi_araddr        ),
  .m23_axi_arlen         ( m23_axi_arlen         ),
  .m23_axi_rvalid        ( m23_axi_rvalid        ),
  .m23_axi_rready        ( m23_axi_rready        ),
  .m23_axi_rdata         ( m23_axi_rdata         ),
  .m23_axi_rlast         ( m23_axi_rlast         ),
  .m24_axi_awvalid       ( m24_axi_awvalid       ),
  .m24_axi_awready       ( m24_axi_awready       ),
  .m24_axi_awaddr        ( m24_axi_awaddr        ),
  .m24_axi_awlen         ( m24_axi_awlen         ),
  .m24_axi_wvalid        ( m24_axi_wvalid        ),
  .m24_axi_wready        ( m24_axi_wready        ),
  .m24_axi_wdata         ( m24_axi_wdata         ),
  .m24_axi_wstrb         ( m24_axi_wstrb         ),
  .m24_axi_wlast         ( m24_axi_wlast         ),
  .m24_axi_bvalid        ( m24_axi_bvalid        ),
  .m24_axi_bready        ( m24_axi_bready        ),
  .m24_axi_arvalid       ( m24_axi_arvalid       ),
  .m24_axi_arready       ( m24_axi_arready       ),
  .m24_axi_araddr        ( m24_axi_araddr        ),
  .m24_axi_arlen         ( m24_axi_arlen         ),
  .m24_axi_rvalid        ( m24_axi_rvalid        ),
  .m24_axi_rready        ( m24_axi_rready        ),
  .m24_axi_rdata         ( m24_axi_rdata         ),
  .m24_axi_rlast         ( m24_axi_rlast         ),
  .m25_axi_awvalid       ( m25_axi_awvalid       ),
  .m25_axi_awready       ( m25_axi_awready       ),
  .m25_axi_awaddr        ( m25_axi_awaddr        ),
  .m25_axi_awlen         ( m25_axi_awlen         ),
  .m25_axi_wvalid        ( m25_axi_wvalid        ),
  .m25_axi_wready        ( m25_axi_wready        ),
  .m25_axi_wdata         ( m25_axi_wdata         ),
  .m25_axi_wstrb         ( m25_axi_wstrb         ),
  .m25_axi_wlast         ( m25_axi_wlast         ),
  .m25_axi_bvalid        ( m25_axi_bvalid        ),
  .m25_axi_bready        ( m25_axi_bready        ),
  .m25_axi_arvalid       ( m25_axi_arvalid       ),
  .m25_axi_arready       ( m25_axi_arready       ),
  .m25_axi_araddr        ( m25_axi_araddr        ),
  .m25_axi_arlen         ( m25_axi_arlen         ),
  .m25_axi_rvalid        ( m25_axi_rvalid        ),
  .m25_axi_rready        ( m25_axi_rready        ),
  .m25_axi_rdata         ( m25_axi_rdata         ),
  .m25_axi_rlast         ( m25_axi_rlast         ),
  .m26_axi_awvalid       ( m26_axi_awvalid       ),
  .m26_axi_awready       ( m26_axi_awready       ),
  .m26_axi_awaddr        ( m26_axi_awaddr        ),
  .m26_axi_awlen         ( m26_axi_awlen         ),
  .m26_axi_wvalid        ( m26_axi_wvalid        ),
  .m26_axi_wready        ( m26_axi_wready        ),
  .m26_axi_wdata         ( m26_axi_wdata         ),
  .m26_axi_wstrb         ( m26_axi_wstrb         ),
  .m26_axi_wlast         ( m26_axi_wlast         ),
  .m26_axi_bvalid        ( m26_axi_bvalid        ),
  .m26_axi_bready        ( m26_axi_bready        ),
  .m26_axi_arvalid       ( m26_axi_arvalid       ),
  .m26_axi_arready       ( m26_axi_arready       ),
  .m26_axi_araddr        ( m26_axi_araddr        ),
  .m26_axi_arlen         ( m26_axi_arlen         ),
  .m26_axi_rvalid        ( m26_axi_rvalid        ),
  .m26_axi_rready        ( m26_axi_rready        ),
  .m26_axi_rdata         ( m26_axi_rdata         ),
  .m26_axi_rlast         ( m26_axi_rlast         ),
  .m27_axi_awvalid       ( m27_axi_awvalid       ),
  .m27_axi_awready       ( m27_axi_awready       ),
  .m27_axi_awaddr        ( m27_axi_awaddr        ),
  .m27_axi_awlen         ( m27_axi_awlen         ),
  .m27_axi_wvalid        ( m27_axi_wvalid        ),
  .m27_axi_wready        ( m27_axi_wready        ),
  .m27_axi_wdata         ( m27_axi_wdata         ),
  .m27_axi_wstrb         ( m27_axi_wstrb         ),
  .m27_axi_wlast         ( m27_axi_wlast         ),
  .m27_axi_bvalid        ( m27_axi_bvalid        ),
  .m27_axi_bready        ( m27_axi_bready        ),
  .m27_axi_arvalid       ( m27_axi_arvalid       ),
  .m27_axi_arready       ( m27_axi_arready       ),
  .m27_axi_araddr        ( m27_axi_araddr        ),
  .m27_axi_arlen         ( m27_axi_arlen         ),
  .m27_axi_rvalid        ( m27_axi_rvalid        ),
  .m27_axi_rready        ( m27_axi_rready        ),
  .m27_axi_rdata         ( m27_axi_rdata         ),
  .m27_axi_rlast         ( m27_axi_rlast         ),
  .m28_axi_awvalid       ( m28_axi_awvalid       ),
  .m28_axi_awready       ( m28_axi_awready       ),
  .m28_axi_awaddr        ( m28_axi_awaddr        ),
  .m28_axi_awlen         ( m28_axi_awlen         ),
  .m28_axi_wvalid        ( m28_axi_wvalid        ),
  .m28_axi_wready        ( m28_axi_wready        ),
  .m28_axi_wdata         ( m28_axi_wdata         ),
  .m28_axi_wstrb         ( m28_axi_wstrb         ),
  .m28_axi_wlast         ( m28_axi_wlast         ),
  .m28_axi_bvalid        ( m28_axi_bvalid        ),
  .m28_axi_bready        ( m28_axi_bready        ),
  .m28_axi_arvalid       ( m28_axi_arvalid       ),
  .m28_axi_arready       ( m28_axi_arready       ),
  .m28_axi_araddr        ( m28_axi_araddr        ),
  .m28_axi_arlen         ( m28_axi_arlen         ),
  .m28_axi_rvalid        ( m28_axi_rvalid        ),
  .m28_axi_rready        ( m28_axi_rready        ),
  .m28_axi_rdata         ( m28_axi_rdata         ),
  .m28_axi_rlast         ( m28_axi_rlast         ),
  .m29_axi_awvalid       ( m29_axi_awvalid       ),
  .m29_axi_awready       ( m29_axi_awready       ),
  .m29_axi_awaddr        ( m29_axi_awaddr        ),
  .m29_axi_awlen         ( m29_axi_awlen         ),
  .m29_axi_wvalid        ( m29_axi_wvalid        ),
  .m29_axi_wready        ( m29_axi_wready        ),
  .m29_axi_wdata         ( m29_axi_wdata         ),
  .m29_axi_wstrb         ( m29_axi_wstrb         ),
  .m29_axi_wlast         ( m29_axi_wlast         ),
  .m29_axi_bvalid        ( m29_axi_bvalid        ),
  .m29_axi_bready        ( m29_axi_bready        ),
  .m29_axi_arvalid       ( m29_axi_arvalid       ),
  .m29_axi_arready       ( m29_axi_arready       ),
  .m29_axi_araddr        ( m29_axi_araddr        ),
  .m29_axi_arlen         ( m29_axi_arlen         ),
  .m29_axi_rvalid        ( m29_axi_rvalid        ),
  .m29_axi_rready        ( m29_axi_rready        ),
  .m29_axi_rdata         ( m29_axi_rdata         ),
  .m29_axi_rlast         ( m29_axi_rlast         ),
  .m30_axi_awvalid       ( m30_axi_awvalid       ),
  .m30_axi_awready       ( m30_axi_awready       ),
  .m30_axi_awaddr        ( m30_axi_awaddr        ),
  .m30_axi_awlen         ( m30_axi_awlen         ),
  .m30_axi_wvalid        ( m30_axi_wvalid        ),
  .m30_axi_wready        ( m30_axi_wready        ),
  .m30_axi_wdata         ( m30_axi_wdata         ),
  .m30_axi_wstrb         ( m30_axi_wstrb         ),
  .m30_axi_wlast         ( m30_axi_wlast         ),
  .m30_axi_bvalid        ( m30_axi_bvalid        ),
  .m30_axi_bready        ( m30_axi_bready        ),
  .m30_axi_arvalid       ( m30_axi_arvalid       ),
  .m30_axi_arready       ( m30_axi_arready       ),
  .m30_axi_araddr        ( m30_axi_araddr        ),
  .m30_axi_arlen         ( m30_axi_arlen         ),
  .m30_axi_rvalid        ( m30_axi_rvalid        ),
  .m30_axi_rready        ( m30_axi_rready        ),
  .m30_axi_rdata         ( m30_axi_rdata         ),
  .m30_axi_rlast         ( m30_axi_rlast         ),
  .m31_axi_awvalid       ( m31_axi_awvalid       ),
  .m31_axi_awready       ( m31_axi_awready       ),
  .m31_axi_awaddr        ( m31_axi_awaddr        ),
  .m31_axi_awlen         ( m31_axi_awlen         ),
  .m31_axi_wvalid        ( m31_axi_wvalid        ),
  .m31_axi_wready        ( m31_axi_wready        ),
  .m31_axi_wdata         ( m31_axi_wdata         ),
  .m31_axi_wstrb         ( m31_axi_wstrb         ),
  .m31_axi_wlast         ( m31_axi_wlast         ),
  .m31_axi_bvalid        ( m31_axi_bvalid        ),
  .m31_axi_bready        ( m31_axi_bready        ),
  .m31_axi_arvalid       ( m31_axi_arvalid       ),
  .m31_axi_arready       ( m31_axi_arready       ),
  .m31_axi_araddr        ( m31_axi_araddr        ),
  .m31_axi_arlen         ( m31_axi_arlen         ),
  .m31_axi_rvalid        ( m31_axi_rvalid        ),
  .m31_axi_rready        ( m31_axi_rready        ),
  .m31_axi_rdata         ( m31_axi_rdata         ),
  .m31_axi_rlast         ( m31_axi_rlast         ),
  .s_axi_control_awvalid ( s_axi_control_awvalid ),
  .s_axi_control_awready ( s_axi_control_awready ),
  .s_axi_control_awaddr  ( s_axi_control_awaddr  ),
  .s_axi_control_wvalid  ( s_axi_control_wvalid  ),
  .s_axi_control_wready  ( s_axi_control_wready  ),
  .s_axi_control_wdata   ( s_axi_control_wdata   ),
  .s_axi_control_wstrb   ( s_axi_control_wstrb   ),
  .s_axi_control_arvalid ( s_axi_control_arvalid ),
  .s_axi_control_arready ( s_axi_control_arready ),
  .s_axi_control_araddr  ( s_axi_control_araddr  ),
  .s_axi_control_rvalid  ( s_axi_control_rvalid  ),
  .s_axi_control_rready  ( s_axi_control_rready  ),
  .s_axi_control_rdata   ( s_axi_control_rdata   ),
  .s_axi_control_rresp   ( s_axi_control_rresp   ),
  .s_axi_control_bvalid  ( s_axi_control_bvalid  ),
  .s_axi_control_bready  ( s_axi_control_bready  ),
  .s_axi_control_bresp   ( s_axi_control_bresp   ),
  .interrupt             ( interrupt             )
);

// Master Control instantiation
control_acc_kernel_vip inst_control_acc_kernel_vip (
  .aclk          ( ap_clk                ),
  .aresetn       ( ap_rst_n              ),
  .m_axi_awvalid ( s_axi_control_awvalid ),
  .m_axi_awready ( s_axi_control_awready ),
  .m_axi_awaddr  ( s_axi_control_awaddr  ),
  .m_axi_wvalid  ( s_axi_control_wvalid  ),
  .m_axi_wready  ( s_axi_control_wready  ),
  .m_axi_wdata   ( s_axi_control_wdata   ),
  .m_axi_wstrb   ( s_axi_control_wstrb   ),
  .m_axi_arvalid ( s_axi_control_arvalid ),
  .m_axi_arready ( s_axi_control_arready ),
  .m_axi_araddr  ( s_axi_control_araddr  ),
  .m_axi_rvalid  ( s_axi_control_rvalid  ),
  .m_axi_rready  ( s_axi_control_rready  ),
  .m_axi_rdata   ( s_axi_control_rdata   ),
  .m_axi_rresp   ( s_axi_control_rresp   ),
  .m_axi_bvalid  ( s_axi_control_bvalid  ),
  .m_axi_bready  ( s_axi_control_bready  ),
  .m_axi_bresp   ( s_axi_control_bresp   )
);

control_acc_kernel_vip_mst_t  ctrl;

// Slave MM VIP instantiation
slv_m00_axi_vip inst_slv_m00_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m00_axi_awvalid ),
  .s_axi_awready ( m00_axi_awready ),
  .s_axi_awaddr  ( m00_axi_awaddr  ),
  .s_axi_awlen   ( m00_axi_awlen   ),
  .s_axi_wvalid  ( m00_axi_wvalid  ),
  .s_axi_wready  ( m00_axi_wready  ),
  .s_axi_wdata   ( m00_axi_wdata   ),
  .s_axi_wstrb   ( m00_axi_wstrb   ),
  .s_axi_wlast   ( m00_axi_wlast   ),
  .s_axi_bvalid  ( m00_axi_bvalid  ),
  .s_axi_bready  ( m00_axi_bready  ),
  .s_axi_arvalid ( m00_axi_arvalid ),
  .s_axi_arready ( m00_axi_arready ),
  .s_axi_araddr  ( m00_axi_araddr  ),
  .s_axi_arlen   ( m00_axi_arlen   ),
  .s_axi_rvalid  ( m00_axi_rvalid  ),
  .s_axi_rready  ( m00_axi_rready  ),
  .s_axi_rdata   ( m00_axi_rdata   ),
  .s_axi_rlast   ( m00_axi_rlast   )
);


slv_m00_axi_vip_slv_mem_t   m00_axi;
slv_m00_axi_vip_slv_t   m00_axi_slv;

// Slave MM VIP instantiation
slv_m01_axi_vip inst_slv_m01_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m01_axi_awvalid ),
  .s_axi_awready ( m01_axi_awready ),
  .s_axi_awaddr  ( m01_axi_awaddr  ),
  .s_axi_awlen   ( m01_axi_awlen   ),
  .s_axi_wvalid  ( m01_axi_wvalid  ),
  .s_axi_wready  ( m01_axi_wready  ),
  .s_axi_wdata   ( m01_axi_wdata   ),
  .s_axi_wstrb   ( m01_axi_wstrb   ),
  .s_axi_wlast   ( m01_axi_wlast   ),
  .s_axi_bvalid  ( m01_axi_bvalid  ),
  .s_axi_bready  ( m01_axi_bready  ),
  .s_axi_arvalid ( m01_axi_arvalid ),
  .s_axi_arready ( m01_axi_arready ),
  .s_axi_araddr  ( m01_axi_araddr  ),
  .s_axi_arlen   ( m01_axi_arlen   ),
  .s_axi_rvalid  ( m01_axi_rvalid  ),
  .s_axi_rready  ( m01_axi_rready  ),
  .s_axi_rdata   ( m01_axi_rdata   ),
  .s_axi_rlast   ( m01_axi_rlast   )
);


slv_m01_axi_vip_slv_mem_t   m01_axi;
slv_m01_axi_vip_slv_t   m01_axi_slv;

// Slave MM VIP instantiation
slv_m02_axi_vip inst_slv_m02_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m02_axi_awvalid ),
  .s_axi_awready ( m02_axi_awready ),
  .s_axi_awaddr  ( m02_axi_awaddr  ),
  .s_axi_awlen   ( m02_axi_awlen   ),
  .s_axi_wvalid  ( m02_axi_wvalid  ),
  .s_axi_wready  ( m02_axi_wready  ),
  .s_axi_wdata   ( m02_axi_wdata   ),
  .s_axi_wstrb   ( m02_axi_wstrb   ),
  .s_axi_wlast   ( m02_axi_wlast   ),
  .s_axi_bvalid  ( m02_axi_bvalid  ),
  .s_axi_bready  ( m02_axi_bready  ),
  .s_axi_arvalid ( m02_axi_arvalid ),
  .s_axi_arready ( m02_axi_arready ),
  .s_axi_araddr  ( m02_axi_araddr  ),
  .s_axi_arlen   ( m02_axi_arlen   ),
  .s_axi_rvalid  ( m02_axi_rvalid  ),
  .s_axi_rready  ( m02_axi_rready  ),
  .s_axi_rdata   ( m02_axi_rdata   ),
  .s_axi_rlast   ( m02_axi_rlast   )
);


slv_m02_axi_vip_slv_mem_t   m02_axi;
slv_m02_axi_vip_slv_t   m02_axi_slv;

// Slave MM VIP instantiation
slv_m03_axi_vip inst_slv_m03_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m03_axi_awvalid ),
  .s_axi_awready ( m03_axi_awready ),
  .s_axi_awaddr  ( m03_axi_awaddr  ),
  .s_axi_awlen   ( m03_axi_awlen   ),
  .s_axi_wvalid  ( m03_axi_wvalid  ),
  .s_axi_wready  ( m03_axi_wready  ),
  .s_axi_wdata   ( m03_axi_wdata   ),
  .s_axi_wstrb   ( m03_axi_wstrb   ),
  .s_axi_wlast   ( m03_axi_wlast   ),
  .s_axi_bvalid  ( m03_axi_bvalid  ),
  .s_axi_bready  ( m03_axi_bready  ),
  .s_axi_arvalid ( m03_axi_arvalid ),
  .s_axi_arready ( m03_axi_arready ),
  .s_axi_araddr  ( m03_axi_araddr  ),
  .s_axi_arlen   ( m03_axi_arlen   ),
  .s_axi_rvalid  ( m03_axi_rvalid  ),
  .s_axi_rready  ( m03_axi_rready  ),
  .s_axi_rdata   ( m03_axi_rdata   ),
  .s_axi_rlast   ( m03_axi_rlast   )
);


slv_m03_axi_vip_slv_mem_t   m03_axi;
slv_m03_axi_vip_slv_t   m03_axi_slv;

// Slave MM VIP instantiation
slv_m04_axi_vip inst_slv_m04_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m04_axi_awvalid ),
  .s_axi_awready ( m04_axi_awready ),
  .s_axi_awaddr  ( m04_axi_awaddr  ),
  .s_axi_awlen   ( m04_axi_awlen   ),
  .s_axi_wvalid  ( m04_axi_wvalid  ),
  .s_axi_wready  ( m04_axi_wready  ),
  .s_axi_wdata   ( m04_axi_wdata   ),
  .s_axi_wstrb   ( m04_axi_wstrb   ),
  .s_axi_wlast   ( m04_axi_wlast   ),
  .s_axi_bvalid  ( m04_axi_bvalid  ),
  .s_axi_bready  ( m04_axi_bready  ),
  .s_axi_arvalid ( m04_axi_arvalid ),
  .s_axi_arready ( m04_axi_arready ),
  .s_axi_araddr  ( m04_axi_araddr  ),
  .s_axi_arlen   ( m04_axi_arlen   ),
  .s_axi_rvalid  ( m04_axi_rvalid  ),
  .s_axi_rready  ( m04_axi_rready  ),
  .s_axi_rdata   ( m04_axi_rdata   ),
  .s_axi_rlast   ( m04_axi_rlast   )
);


slv_m04_axi_vip_slv_mem_t   m04_axi;
slv_m04_axi_vip_slv_t   m04_axi_slv;

// Slave MM VIP instantiation
slv_m05_axi_vip inst_slv_m05_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m05_axi_awvalid ),
  .s_axi_awready ( m05_axi_awready ),
  .s_axi_awaddr  ( m05_axi_awaddr  ),
  .s_axi_awlen   ( m05_axi_awlen   ),
  .s_axi_wvalid  ( m05_axi_wvalid  ),
  .s_axi_wready  ( m05_axi_wready  ),
  .s_axi_wdata   ( m05_axi_wdata   ),
  .s_axi_wstrb   ( m05_axi_wstrb   ),
  .s_axi_wlast   ( m05_axi_wlast   ),
  .s_axi_bvalid  ( m05_axi_bvalid  ),
  .s_axi_bready  ( m05_axi_bready  ),
  .s_axi_arvalid ( m05_axi_arvalid ),
  .s_axi_arready ( m05_axi_arready ),
  .s_axi_araddr  ( m05_axi_araddr  ),
  .s_axi_arlen   ( m05_axi_arlen   ),
  .s_axi_rvalid  ( m05_axi_rvalid  ),
  .s_axi_rready  ( m05_axi_rready  ),
  .s_axi_rdata   ( m05_axi_rdata   ),
  .s_axi_rlast   ( m05_axi_rlast   )
);


slv_m05_axi_vip_slv_mem_t   m05_axi;
slv_m05_axi_vip_slv_t   m05_axi_slv;

// Slave MM VIP instantiation
slv_m06_axi_vip inst_slv_m06_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m06_axi_awvalid ),
  .s_axi_awready ( m06_axi_awready ),
  .s_axi_awaddr  ( m06_axi_awaddr  ),
  .s_axi_awlen   ( m06_axi_awlen   ),
  .s_axi_wvalid  ( m06_axi_wvalid  ),
  .s_axi_wready  ( m06_axi_wready  ),
  .s_axi_wdata   ( m06_axi_wdata   ),
  .s_axi_wstrb   ( m06_axi_wstrb   ),
  .s_axi_wlast   ( m06_axi_wlast   ),
  .s_axi_bvalid  ( m06_axi_bvalid  ),
  .s_axi_bready  ( m06_axi_bready  ),
  .s_axi_arvalid ( m06_axi_arvalid ),
  .s_axi_arready ( m06_axi_arready ),
  .s_axi_araddr  ( m06_axi_araddr  ),
  .s_axi_arlen   ( m06_axi_arlen   ),
  .s_axi_rvalid  ( m06_axi_rvalid  ),
  .s_axi_rready  ( m06_axi_rready  ),
  .s_axi_rdata   ( m06_axi_rdata   ),
  .s_axi_rlast   ( m06_axi_rlast   )
);


slv_m06_axi_vip_slv_mem_t   m06_axi;
slv_m06_axi_vip_slv_t   m06_axi_slv;

// Slave MM VIP instantiation
slv_m07_axi_vip inst_slv_m07_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m07_axi_awvalid ),
  .s_axi_awready ( m07_axi_awready ),
  .s_axi_awaddr  ( m07_axi_awaddr  ),
  .s_axi_awlen   ( m07_axi_awlen   ),
  .s_axi_wvalid  ( m07_axi_wvalid  ),
  .s_axi_wready  ( m07_axi_wready  ),
  .s_axi_wdata   ( m07_axi_wdata   ),
  .s_axi_wstrb   ( m07_axi_wstrb   ),
  .s_axi_wlast   ( m07_axi_wlast   ),
  .s_axi_bvalid  ( m07_axi_bvalid  ),
  .s_axi_bready  ( m07_axi_bready  ),
  .s_axi_arvalid ( m07_axi_arvalid ),
  .s_axi_arready ( m07_axi_arready ),
  .s_axi_araddr  ( m07_axi_araddr  ),
  .s_axi_arlen   ( m07_axi_arlen   ),
  .s_axi_rvalid  ( m07_axi_rvalid  ),
  .s_axi_rready  ( m07_axi_rready  ),
  .s_axi_rdata   ( m07_axi_rdata   ),
  .s_axi_rlast   ( m07_axi_rlast   )
);


slv_m07_axi_vip_slv_mem_t   m07_axi;
slv_m07_axi_vip_slv_t   m07_axi_slv;

// Slave MM VIP instantiation
slv_m08_axi_vip inst_slv_m08_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m08_axi_awvalid ),
  .s_axi_awready ( m08_axi_awready ),
  .s_axi_awaddr  ( m08_axi_awaddr  ),
  .s_axi_awlen   ( m08_axi_awlen   ),
  .s_axi_wvalid  ( m08_axi_wvalid  ),
  .s_axi_wready  ( m08_axi_wready  ),
  .s_axi_wdata   ( m08_axi_wdata   ),
  .s_axi_wstrb   ( m08_axi_wstrb   ),
  .s_axi_wlast   ( m08_axi_wlast   ),
  .s_axi_bvalid  ( m08_axi_bvalid  ),
  .s_axi_bready  ( m08_axi_bready  ),
  .s_axi_arvalid ( m08_axi_arvalid ),
  .s_axi_arready ( m08_axi_arready ),
  .s_axi_araddr  ( m08_axi_araddr  ),
  .s_axi_arlen   ( m08_axi_arlen   ),
  .s_axi_rvalid  ( m08_axi_rvalid  ),
  .s_axi_rready  ( m08_axi_rready  ),
  .s_axi_rdata   ( m08_axi_rdata   ),
  .s_axi_rlast   ( m08_axi_rlast   )
);


slv_m08_axi_vip_slv_mem_t   m08_axi;
slv_m08_axi_vip_slv_t   m08_axi_slv;

// Slave MM VIP instantiation
slv_m09_axi_vip inst_slv_m09_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m09_axi_awvalid ),
  .s_axi_awready ( m09_axi_awready ),
  .s_axi_awaddr  ( m09_axi_awaddr  ),
  .s_axi_awlen   ( m09_axi_awlen   ),
  .s_axi_wvalid  ( m09_axi_wvalid  ),
  .s_axi_wready  ( m09_axi_wready  ),
  .s_axi_wdata   ( m09_axi_wdata   ),
  .s_axi_wstrb   ( m09_axi_wstrb   ),
  .s_axi_wlast   ( m09_axi_wlast   ),
  .s_axi_bvalid  ( m09_axi_bvalid  ),
  .s_axi_bready  ( m09_axi_bready  ),
  .s_axi_arvalid ( m09_axi_arvalid ),
  .s_axi_arready ( m09_axi_arready ),
  .s_axi_araddr  ( m09_axi_araddr  ),
  .s_axi_arlen   ( m09_axi_arlen   ),
  .s_axi_rvalid  ( m09_axi_rvalid  ),
  .s_axi_rready  ( m09_axi_rready  ),
  .s_axi_rdata   ( m09_axi_rdata   ),
  .s_axi_rlast   ( m09_axi_rlast   )
);


slv_m09_axi_vip_slv_mem_t   m09_axi;
slv_m09_axi_vip_slv_t   m09_axi_slv;

// Slave MM VIP instantiation
slv_m10_axi_vip inst_slv_m10_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m10_axi_awvalid ),
  .s_axi_awready ( m10_axi_awready ),
  .s_axi_awaddr  ( m10_axi_awaddr  ),
  .s_axi_awlen   ( m10_axi_awlen   ),
  .s_axi_wvalid  ( m10_axi_wvalid  ),
  .s_axi_wready  ( m10_axi_wready  ),
  .s_axi_wdata   ( m10_axi_wdata   ),
  .s_axi_wstrb   ( m10_axi_wstrb   ),
  .s_axi_wlast   ( m10_axi_wlast   ),
  .s_axi_bvalid  ( m10_axi_bvalid  ),
  .s_axi_bready  ( m10_axi_bready  ),
  .s_axi_arvalid ( m10_axi_arvalid ),
  .s_axi_arready ( m10_axi_arready ),
  .s_axi_araddr  ( m10_axi_araddr  ),
  .s_axi_arlen   ( m10_axi_arlen   ),
  .s_axi_rvalid  ( m10_axi_rvalid  ),
  .s_axi_rready  ( m10_axi_rready  ),
  .s_axi_rdata   ( m10_axi_rdata   ),
  .s_axi_rlast   ( m10_axi_rlast   )
);


slv_m10_axi_vip_slv_mem_t   m10_axi;
slv_m10_axi_vip_slv_t   m10_axi_slv;

// Slave MM VIP instantiation
slv_m11_axi_vip inst_slv_m11_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m11_axi_awvalid ),
  .s_axi_awready ( m11_axi_awready ),
  .s_axi_awaddr  ( m11_axi_awaddr  ),
  .s_axi_awlen   ( m11_axi_awlen   ),
  .s_axi_wvalid  ( m11_axi_wvalid  ),
  .s_axi_wready  ( m11_axi_wready  ),
  .s_axi_wdata   ( m11_axi_wdata   ),
  .s_axi_wstrb   ( m11_axi_wstrb   ),
  .s_axi_wlast   ( m11_axi_wlast   ),
  .s_axi_bvalid  ( m11_axi_bvalid  ),
  .s_axi_bready  ( m11_axi_bready  ),
  .s_axi_arvalid ( m11_axi_arvalid ),
  .s_axi_arready ( m11_axi_arready ),
  .s_axi_araddr  ( m11_axi_araddr  ),
  .s_axi_arlen   ( m11_axi_arlen   ),
  .s_axi_rvalid  ( m11_axi_rvalid  ),
  .s_axi_rready  ( m11_axi_rready  ),
  .s_axi_rdata   ( m11_axi_rdata   ),
  .s_axi_rlast   ( m11_axi_rlast   )
);


slv_m11_axi_vip_slv_mem_t   m11_axi;
slv_m11_axi_vip_slv_t   m11_axi_slv;

// Slave MM VIP instantiation
slv_m12_axi_vip inst_slv_m12_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m12_axi_awvalid ),
  .s_axi_awready ( m12_axi_awready ),
  .s_axi_awaddr  ( m12_axi_awaddr  ),
  .s_axi_awlen   ( m12_axi_awlen   ),
  .s_axi_wvalid  ( m12_axi_wvalid  ),
  .s_axi_wready  ( m12_axi_wready  ),
  .s_axi_wdata   ( m12_axi_wdata   ),
  .s_axi_wstrb   ( m12_axi_wstrb   ),
  .s_axi_wlast   ( m12_axi_wlast   ),
  .s_axi_bvalid  ( m12_axi_bvalid  ),
  .s_axi_bready  ( m12_axi_bready  ),
  .s_axi_arvalid ( m12_axi_arvalid ),
  .s_axi_arready ( m12_axi_arready ),
  .s_axi_araddr  ( m12_axi_araddr  ),
  .s_axi_arlen   ( m12_axi_arlen   ),
  .s_axi_rvalid  ( m12_axi_rvalid  ),
  .s_axi_rready  ( m12_axi_rready  ),
  .s_axi_rdata   ( m12_axi_rdata   ),
  .s_axi_rlast   ( m12_axi_rlast   )
);


slv_m12_axi_vip_slv_mem_t   m12_axi;
slv_m12_axi_vip_slv_t   m12_axi_slv;

// Slave MM VIP instantiation
slv_m13_axi_vip inst_slv_m13_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m13_axi_awvalid ),
  .s_axi_awready ( m13_axi_awready ),
  .s_axi_awaddr  ( m13_axi_awaddr  ),
  .s_axi_awlen   ( m13_axi_awlen   ),
  .s_axi_wvalid  ( m13_axi_wvalid  ),
  .s_axi_wready  ( m13_axi_wready  ),
  .s_axi_wdata   ( m13_axi_wdata   ),
  .s_axi_wstrb   ( m13_axi_wstrb   ),
  .s_axi_wlast   ( m13_axi_wlast   ),
  .s_axi_bvalid  ( m13_axi_bvalid  ),
  .s_axi_bready  ( m13_axi_bready  ),
  .s_axi_arvalid ( m13_axi_arvalid ),
  .s_axi_arready ( m13_axi_arready ),
  .s_axi_araddr  ( m13_axi_araddr  ),
  .s_axi_arlen   ( m13_axi_arlen   ),
  .s_axi_rvalid  ( m13_axi_rvalid  ),
  .s_axi_rready  ( m13_axi_rready  ),
  .s_axi_rdata   ( m13_axi_rdata   ),
  .s_axi_rlast   ( m13_axi_rlast   )
);


slv_m13_axi_vip_slv_mem_t   m13_axi;
slv_m13_axi_vip_slv_t   m13_axi_slv;

// Slave MM VIP instantiation
slv_m14_axi_vip inst_slv_m14_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m14_axi_awvalid ),
  .s_axi_awready ( m14_axi_awready ),
  .s_axi_awaddr  ( m14_axi_awaddr  ),
  .s_axi_awlen   ( m14_axi_awlen   ),
  .s_axi_wvalid  ( m14_axi_wvalid  ),
  .s_axi_wready  ( m14_axi_wready  ),
  .s_axi_wdata   ( m14_axi_wdata   ),
  .s_axi_wstrb   ( m14_axi_wstrb   ),
  .s_axi_wlast   ( m14_axi_wlast   ),
  .s_axi_bvalid  ( m14_axi_bvalid  ),
  .s_axi_bready  ( m14_axi_bready  ),
  .s_axi_arvalid ( m14_axi_arvalid ),
  .s_axi_arready ( m14_axi_arready ),
  .s_axi_araddr  ( m14_axi_araddr  ),
  .s_axi_arlen   ( m14_axi_arlen   ),
  .s_axi_rvalid  ( m14_axi_rvalid  ),
  .s_axi_rready  ( m14_axi_rready  ),
  .s_axi_rdata   ( m14_axi_rdata   ),
  .s_axi_rlast   ( m14_axi_rlast   )
);


slv_m14_axi_vip_slv_mem_t   m14_axi;
slv_m14_axi_vip_slv_t   m14_axi_slv;

// Slave MM VIP instantiation
slv_m15_axi_vip inst_slv_m15_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m15_axi_awvalid ),
  .s_axi_awready ( m15_axi_awready ),
  .s_axi_awaddr  ( m15_axi_awaddr  ),
  .s_axi_awlen   ( m15_axi_awlen   ),
  .s_axi_wvalid  ( m15_axi_wvalid  ),
  .s_axi_wready  ( m15_axi_wready  ),
  .s_axi_wdata   ( m15_axi_wdata   ),
  .s_axi_wstrb   ( m15_axi_wstrb   ),
  .s_axi_wlast   ( m15_axi_wlast   ),
  .s_axi_bvalid  ( m15_axi_bvalid  ),
  .s_axi_bready  ( m15_axi_bready  ),
  .s_axi_arvalid ( m15_axi_arvalid ),
  .s_axi_arready ( m15_axi_arready ),
  .s_axi_araddr  ( m15_axi_araddr  ),
  .s_axi_arlen   ( m15_axi_arlen   ),
  .s_axi_rvalid  ( m15_axi_rvalid  ),
  .s_axi_rready  ( m15_axi_rready  ),
  .s_axi_rdata   ( m15_axi_rdata   ),
  .s_axi_rlast   ( m15_axi_rlast   )
);


slv_m15_axi_vip_slv_mem_t   m15_axi;
slv_m15_axi_vip_slv_t   m15_axi_slv;

// Slave MM VIP instantiation
slv_m16_axi_vip inst_slv_m16_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m16_axi_awvalid ),
  .s_axi_awready ( m16_axi_awready ),
  .s_axi_awaddr  ( m16_axi_awaddr  ),
  .s_axi_awlen   ( m16_axi_awlen   ),
  .s_axi_wvalid  ( m16_axi_wvalid  ),
  .s_axi_wready  ( m16_axi_wready  ),
  .s_axi_wdata   ( m16_axi_wdata   ),
  .s_axi_wstrb   ( m16_axi_wstrb   ),
  .s_axi_wlast   ( m16_axi_wlast   ),
  .s_axi_bvalid  ( m16_axi_bvalid  ),
  .s_axi_bready  ( m16_axi_bready  ),
  .s_axi_arvalid ( m16_axi_arvalid ),
  .s_axi_arready ( m16_axi_arready ),
  .s_axi_araddr  ( m16_axi_araddr  ),
  .s_axi_arlen   ( m16_axi_arlen   ),
  .s_axi_rvalid  ( m16_axi_rvalid  ),
  .s_axi_rready  ( m16_axi_rready  ),
  .s_axi_rdata   ( m16_axi_rdata   ),
  .s_axi_rlast   ( m16_axi_rlast   )
);


slv_m16_axi_vip_slv_mem_t   m16_axi;
slv_m16_axi_vip_slv_t   m16_axi_slv;

// Slave MM VIP instantiation
slv_m17_axi_vip inst_slv_m17_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m17_axi_awvalid ),
  .s_axi_awready ( m17_axi_awready ),
  .s_axi_awaddr  ( m17_axi_awaddr  ),
  .s_axi_awlen   ( m17_axi_awlen   ),
  .s_axi_wvalid  ( m17_axi_wvalid  ),
  .s_axi_wready  ( m17_axi_wready  ),
  .s_axi_wdata   ( m17_axi_wdata   ),
  .s_axi_wstrb   ( m17_axi_wstrb   ),
  .s_axi_wlast   ( m17_axi_wlast   ),
  .s_axi_bvalid  ( m17_axi_bvalid  ),
  .s_axi_bready  ( m17_axi_bready  ),
  .s_axi_arvalid ( m17_axi_arvalid ),
  .s_axi_arready ( m17_axi_arready ),
  .s_axi_araddr  ( m17_axi_araddr  ),
  .s_axi_arlen   ( m17_axi_arlen   ),
  .s_axi_rvalid  ( m17_axi_rvalid  ),
  .s_axi_rready  ( m17_axi_rready  ),
  .s_axi_rdata   ( m17_axi_rdata   ),
  .s_axi_rlast   ( m17_axi_rlast   )
);


slv_m17_axi_vip_slv_mem_t   m17_axi;
slv_m17_axi_vip_slv_t   m17_axi_slv;

// Slave MM VIP instantiation
slv_m18_axi_vip inst_slv_m18_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m18_axi_awvalid ),
  .s_axi_awready ( m18_axi_awready ),
  .s_axi_awaddr  ( m18_axi_awaddr  ),
  .s_axi_awlen   ( m18_axi_awlen   ),
  .s_axi_wvalid  ( m18_axi_wvalid  ),
  .s_axi_wready  ( m18_axi_wready  ),
  .s_axi_wdata   ( m18_axi_wdata   ),
  .s_axi_wstrb   ( m18_axi_wstrb   ),
  .s_axi_wlast   ( m18_axi_wlast   ),
  .s_axi_bvalid  ( m18_axi_bvalid  ),
  .s_axi_bready  ( m18_axi_bready  ),
  .s_axi_arvalid ( m18_axi_arvalid ),
  .s_axi_arready ( m18_axi_arready ),
  .s_axi_araddr  ( m18_axi_araddr  ),
  .s_axi_arlen   ( m18_axi_arlen   ),
  .s_axi_rvalid  ( m18_axi_rvalid  ),
  .s_axi_rready  ( m18_axi_rready  ),
  .s_axi_rdata   ( m18_axi_rdata   ),
  .s_axi_rlast   ( m18_axi_rlast   )
);


slv_m18_axi_vip_slv_mem_t   m18_axi;
slv_m18_axi_vip_slv_t   m18_axi_slv;

// Slave MM VIP instantiation
slv_m19_axi_vip inst_slv_m19_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m19_axi_awvalid ),
  .s_axi_awready ( m19_axi_awready ),
  .s_axi_awaddr  ( m19_axi_awaddr  ),
  .s_axi_awlen   ( m19_axi_awlen   ),
  .s_axi_wvalid  ( m19_axi_wvalid  ),
  .s_axi_wready  ( m19_axi_wready  ),
  .s_axi_wdata   ( m19_axi_wdata   ),
  .s_axi_wstrb   ( m19_axi_wstrb   ),
  .s_axi_wlast   ( m19_axi_wlast   ),
  .s_axi_bvalid  ( m19_axi_bvalid  ),
  .s_axi_bready  ( m19_axi_bready  ),
  .s_axi_arvalid ( m19_axi_arvalid ),
  .s_axi_arready ( m19_axi_arready ),
  .s_axi_araddr  ( m19_axi_araddr  ),
  .s_axi_arlen   ( m19_axi_arlen   ),
  .s_axi_rvalid  ( m19_axi_rvalid  ),
  .s_axi_rready  ( m19_axi_rready  ),
  .s_axi_rdata   ( m19_axi_rdata   ),
  .s_axi_rlast   ( m19_axi_rlast   )
);


slv_m19_axi_vip_slv_mem_t   m19_axi;
slv_m19_axi_vip_slv_t   m19_axi_slv;

// Slave MM VIP instantiation
slv_m20_axi_vip inst_slv_m20_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m20_axi_awvalid ),
  .s_axi_awready ( m20_axi_awready ),
  .s_axi_awaddr  ( m20_axi_awaddr  ),
  .s_axi_awlen   ( m20_axi_awlen   ),
  .s_axi_wvalid  ( m20_axi_wvalid  ),
  .s_axi_wready  ( m20_axi_wready  ),
  .s_axi_wdata   ( m20_axi_wdata   ),
  .s_axi_wstrb   ( m20_axi_wstrb   ),
  .s_axi_wlast   ( m20_axi_wlast   ),
  .s_axi_bvalid  ( m20_axi_bvalid  ),
  .s_axi_bready  ( m20_axi_bready  ),
  .s_axi_arvalid ( m20_axi_arvalid ),
  .s_axi_arready ( m20_axi_arready ),
  .s_axi_araddr  ( m20_axi_araddr  ),
  .s_axi_arlen   ( m20_axi_arlen   ),
  .s_axi_rvalid  ( m20_axi_rvalid  ),
  .s_axi_rready  ( m20_axi_rready  ),
  .s_axi_rdata   ( m20_axi_rdata   ),
  .s_axi_rlast   ( m20_axi_rlast   )
);


slv_m20_axi_vip_slv_mem_t   m20_axi;
slv_m20_axi_vip_slv_t   m20_axi_slv;

// Slave MM VIP instantiation
slv_m21_axi_vip inst_slv_m21_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m21_axi_awvalid ),
  .s_axi_awready ( m21_axi_awready ),
  .s_axi_awaddr  ( m21_axi_awaddr  ),
  .s_axi_awlen   ( m21_axi_awlen   ),
  .s_axi_wvalid  ( m21_axi_wvalid  ),
  .s_axi_wready  ( m21_axi_wready  ),
  .s_axi_wdata   ( m21_axi_wdata   ),
  .s_axi_wstrb   ( m21_axi_wstrb   ),
  .s_axi_wlast   ( m21_axi_wlast   ),
  .s_axi_bvalid  ( m21_axi_bvalid  ),
  .s_axi_bready  ( m21_axi_bready  ),
  .s_axi_arvalid ( m21_axi_arvalid ),
  .s_axi_arready ( m21_axi_arready ),
  .s_axi_araddr  ( m21_axi_araddr  ),
  .s_axi_arlen   ( m21_axi_arlen   ),
  .s_axi_rvalid  ( m21_axi_rvalid  ),
  .s_axi_rready  ( m21_axi_rready  ),
  .s_axi_rdata   ( m21_axi_rdata   ),
  .s_axi_rlast   ( m21_axi_rlast   )
);


slv_m21_axi_vip_slv_mem_t   m21_axi;
slv_m21_axi_vip_slv_t   m21_axi_slv;

// Slave MM VIP instantiation
slv_m22_axi_vip inst_slv_m22_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m22_axi_awvalid ),
  .s_axi_awready ( m22_axi_awready ),
  .s_axi_awaddr  ( m22_axi_awaddr  ),
  .s_axi_awlen   ( m22_axi_awlen   ),
  .s_axi_wvalid  ( m22_axi_wvalid  ),
  .s_axi_wready  ( m22_axi_wready  ),
  .s_axi_wdata   ( m22_axi_wdata   ),
  .s_axi_wstrb   ( m22_axi_wstrb   ),
  .s_axi_wlast   ( m22_axi_wlast   ),
  .s_axi_bvalid  ( m22_axi_bvalid  ),
  .s_axi_bready  ( m22_axi_bready  ),
  .s_axi_arvalid ( m22_axi_arvalid ),
  .s_axi_arready ( m22_axi_arready ),
  .s_axi_araddr  ( m22_axi_araddr  ),
  .s_axi_arlen   ( m22_axi_arlen   ),
  .s_axi_rvalid  ( m22_axi_rvalid  ),
  .s_axi_rready  ( m22_axi_rready  ),
  .s_axi_rdata   ( m22_axi_rdata   ),
  .s_axi_rlast   ( m22_axi_rlast   )
);


slv_m22_axi_vip_slv_mem_t   m22_axi;
slv_m22_axi_vip_slv_t   m22_axi_slv;

// Slave MM VIP instantiation
slv_m23_axi_vip inst_slv_m23_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m23_axi_awvalid ),
  .s_axi_awready ( m23_axi_awready ),
  .s_axi_awaddr  ( m23_axi_awaddr  ),
  .s_axi_awlen   ( m23_axi_awlen   ),
  .s_axi_wvalid  ( m23_axi_wvalid  ),
  .s_axi_wready  ( m23_axi_wready  ),
  .s_axi_wdata   ( m23_axi_wdata   ),
  .s_axi_wstrb   ( m23_axi_wstrb   ),
  .s_axi_wlast   ( m23_axi_wlast   ),
  .s_axi_bvalid  ( m23_axi_bvalid  ),
  .s_axi_bready  ( m23_axi_bready  ),
  .s_axi_arvalid ( m23_axi_arvalid ),
  .s_axi_arready ( m23_axi_arready ),
  .s_axi_araddr  ( m23_axi_araddr  ),
  .s_axi_arlen   ( m23_axi_arlen   ),
  .s_axi_rvalid  ( m23_axi_rvalid  ),
  .s_axi_rready  ( m23_axi_rready  ),
  .s_axi_rdata   ( m23_axi_rdata   ),
  .s_axi_rlast   ( m23_axi_rlast   )
);


slv_m23_axi_vip_slv_mem_t   m23_axi;
slv_m23_axi_vip_slv_t   m23_axi_slv;

// Slave MM VIP instantiation
slv_m24_axi_vip inst_slv_m24_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m24_axi_awvalid ),
  .s_axi_awready ( m24_axi_awready ),
  .s_axi_awaddr  ( m24_axi_awaddr  ),
  .s_axi_awlen   ( m24_axi_awlen   ),
  .s_axi_wvalid  ( m24_axi_wvalid  ),
  .s_axi_wready  ( m24_axi_wready  ),
  .s_axi_wdata   ( m24_axi_wdata   ),
  .s_axi_wstrb   ( m24_axi_wstrb   ),
  .s_axi_wlast   ( m24_axi_wlast   ),
  .s_axi_bvalid  ( m24_axi_bvalid  ),
  .s_axi_bready  ( m24_axi_bready  ),
  .s_axi_arvalid ( m24_axi_arvalid ),
  .s_axi_arready ( m24_axi_arready ),
  .s_axi_araddr  ( m24_axi_araddr  ),
  .s_axi_arlen   ( m24_axi_arlen   ),
  .s_axi_rvalid  ( m24_axi_rvalid  ),
  .s_axi_rready  ( m24_axi_rready  ),
  .s_axi_rdata   ( m24_axi_rdata   ),
  .s_axi_rlast   ( m24_axi_rlast   )
);


slv_m24_axi_vip_slv_mem_t   m24_axi;
slv_m24_axi_vip_slv_t   m24_axi_slv;

// Slave MM VIP instantiation
slv_m25_axi_vip inst_slv_m25_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m25_axi_awvalid ),
  .s_axi_awready ( m25_axi_awready ),
  .s_axi_awaddr  ( m25_axi_awaddr  ),
  .s_axi_awlen   ( m25_axi_awlen   ),
  .s_axi_wvalid  ( m25_axi_wvalid  ),
  .s_axi_wready  ( m25_axi_wready  ),
  .s_axi_wdata   ( m25_axi_wdata   ),
  .s_axi_wstrb   ( m25_axi_wstrb   ),
  .s_axi_wlast   ( m25_axi_wlast   ),
  .s_axi_bvalid  ( m25_axi_bvalid  ),
  .s_axi_bready  ( m25_axi_bready  ),
  .s_axi_arvalid ( m25_axi_arvalid ),
  .s_axi_arready ( m25_axi_arready ),
  .s_axi_araddr  ( m25_axi_araddr  ),
  .s_axi_arlen   ( m25_axi_arlen   ),
  .s_axi_rvalid  ( m25_axi_rvalid  ),
  .s_axi_rready  ( m25_axi_rready  ),
  .s_axi_rdata   ( m25_axi_rdata   ),
  .s_axi_rlast   ( m25_axi_rlast   )
);


slv_m25_axi_vip_slv_mem_t   m25_axi;
slv_m25_axi_vip_slv_t   m25_axi_slv;

// Slave MM VIP instantiation
slv_m26_axi_vip inst_slv_m26_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m26_axi_awvalid ),
  .s_axi_awready ( m26_axi_awready ),
  .s_axi_awaddr  ( m26_axi_awaddr  ),
  .s_axi_awlen   ( m26_axi_awlen   ),
  .s_axi_wvalid  ( m26_axi_wvalid  ),
  .s_axi_wready  ( m26_axi_wready  ),
  .s_axi_wdata   ( m26_axi_wdata   ),
  .s_axi_wstrb   ( m26_axi_wstrb   ),
  .s_axi_wlast   ( m26_axi_wlast   ),
  .s_axi_bvalid  ( m26_axi_bvalid  ),
  .s_axi_bready  ( m26_axi_bready  ),
  .s_axi_arvalid ( m26_axi_arvalid ),
  .s_axi_arready ( m26_axi_arready ),
  .s_axi_araddr  ( m26_axi_araddr  ),
  .s_axi_arlen   ( m26_axi_arlen   ),
  .s_axi_rvalid  ( m26_axi_rvalid  ),
  .s_axi_rready  ( m26_axi_rready  ),
  .s_axi_rdata   ( m26_axi_rdata   ),
  .s_axi_rlast   ( m26_axi_rlast   )
);


slv_m26_axi_vip_slv_mem_t   m26_axi;
slv_m26_axi_vip_slv_t   m26_axi_slv;

// Slave MM VIP instantiation
slv_m27_axi_vip inst_slv_m27_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m27_axi_awvalid ),
  .s_axi_awready ( m27_axi_awready ),
  .s_axi_awaddr  ( m27_axi_awaddr  ),
  .s_axi_awlen   ( m27_axi_awlen   ),
  .s_axi_wvalid  ( m27_axi_wvalid  ),
  .s_axi_wready  ( m27_axi_wready  ),
  .s_axi_wdata   ( m27_axi_wdata   ),
  .s_axi_wstrb   ( m27_axi_wstrb   ),
  .s_axi_wlast   ( m27_axi_wlast   ),
  .s_axi_bvalid  ( m27_axi_bvalid  ),
  .s_axi_bready  ( m27_axi_bready  ),
  .s_axi_arvalid ( m27_axi_arvalid ),
  .s_axi_arready ( m27_axi_arready ),
  .s_axi_araddr  ( m27_axi_araddr  ),
  .s_axi_arlen   ( m27_axi_arlen   ),
  .s_axi_rvalid  ( m27_axi_rvalid  ),
  .s_axi_rready  ( m27_axi_rready  ),
  .s_axi_rdata   ( m27_axi_rdata   ),
  .s_axi_rlast   ( m27_axi_rlast   )
);


slv_m27_axi_vip_slv_mem_t   m27_axi;
slv_m27_axi_vip_slv_t   m27_axi_slv;

// Slave MM VIP instantiation
slv_m28_axi_vip inst_slv_m28_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m28_axi_awvalid ),
  .s_axi_awready ( m28_axi_awready ),
  .s_axi_awaddr  ( m28_axi_awaddr  ),
  .s_axi_awlen   ( m28_axi_awlen   ),
  .s_axi_wvalid  ( m28_axi_wvalid  ),
  .s_axi_wready  ( m28_axi_wready  ),
  .s_axi_wdata   ( m28_axi_wdata   ),
  .s_axi_wstrb   ( m28_axi_wstrb   ),
  .s_axi_wlast   ( m28_axi_wlast   ),
  .s_axi_bvalid  ( m28_axi_bvalid  ),
  .s_axi_bready  ( m28_axi_bready  ),
  .s_axi_arvalid ( m28_axi_arvalid ),
  .s_axi_arready ( m28_axi_arready ),
  .s_axi_araddr  ( m28_axi_araddr  ),
  .s_axi_arlen   ( m28_axi_arlen   ),
  .s_axi_rvalid  ( m28_axi_rvalid  ),
  .s_axi_rready  ( m28_axi_rready  ),
  .s_axi_rdata   ( m28_axi_rdata   ),
  .s_axi_rlast   ( m28_axi_rlast   )
);


slv_m28_axi_vip_slv_mem_t   m28_axi;
slv_m28_axi_vip_slv_t   m28_axi_slv;

// Slave MM VIP instantiation
slv_m29_axi_vip inst_slv_m29_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m29_axi_awvalid ),
  .s_axi_awready ( m29_axi_awready ),
  .s_axi_awaddr  ( m29_axi_awaddr  ),
  .s_axi_awlen   ( m29_axi_awlen   ),
  .s_axi_wvalid  ( m29_axi_wvalid  ),
  .s_axi_wready  ( m29_axi_wready  ),
  .s_axi_wdata   ( m29_axi_wdata   ),
  .s_axi_wstrb   ( m29_axi_wstrb   ),
  .s_axi_wlast   ( m29_axi_wlast   ),
  .s_axi_bvalid  ( m29_axi_bvalid  ),
  .s_axi_bready  ( m29_axi_bready  ),
  .s_axi_arvalid ( m29_axi_arvalid ),
  .s_axi_arready ( m29_axi_arready ),
  .s_axi_araddr  ( m29_axi_araddr  ),
  .s_axi_arlen   ( m29_axi_arlen   ),
  .s_axi_rvalid  ( m29_axi_rvalid  ),
  .s_axi_rready  ( m29_axi_rready  ),
  .s_axi_rdata   ( m29_axi_rdata   ),
  .s_axi_rlast   ( m29_axi_rlast   )
);


slv_m29_axi_vip_slv_mem_t   m29_axi;
slv_m29_axi_vip_slv_t   m29_axi_slv;

// Slave MM VIP instantiation
slv_m30_axi_vip inst_slv_m30_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m30_axi_awvalid ),
  .s_axi_awready ( m30_axi_awready ),
  .s_axi_awaddr  ( m30_axi_awaddr  ),
  .s_axi_awlen   ( m30_axi_awlen   ),
  .s_axi_wvalid  ( m30_axi_wvalid  ),
  .s_axi_wready  ( m30_axi_wready  ),
  .s_axi_wdata   ( m30_axi_wdata   ),
  .s_axi_wstrb   ( m30_axi_wstrb   ),
  .s_axi_wlast   ( m30_axi_wlast   ),
  .s_axi_bvalid  ( m30_axi_bvalid  ),
  .s_axi_bready  ( m30_axi_bready  ),
  .s_axi_arvalid ( m30_axi_arvalid ),
  .s_axi_arready ( m30_axi_arready ),
  .s_axi_araddr  ( m30_axi_araddr  ),
  .s_axi_arlen   ( m30_axi_arlen   ),
  .s_axi_rvalid  ( m30_axi_rvalid  ),
  .s_axi_rready  ( m30_axi_rready  ),
  .s_axi_rdata   ( m30_axi_rdata   ),
  .s_axi_rlast   ( m30_axi_rlast   )
);


slv_m30_axi_vip_slv_mem_t   m30_axi;
slv_m30_axi_vip_slv_t   m30_axi_slv;

// Slave MM VIP instantiation
slv_m31_axi_vip inst_slv_m31_axi_vip (
  .aclk          ( ap_clk          ),
  .aresetn       ( ap_rst_n        ),
  .s_axi_awvalid ( m31_axi_awvalid ),
  .s_axi_awready ( m31_axi_awready ),
  .s_axi_awaddr  ( m31_axi_awaddr  ),
  .s_axi_awlen   ( m31_axi_awlen   ),
  .s_axi_wvalid  ( m31_axi_wvalid  ),
  .s_axi_wready  ( m31_axi_wready  ),
  .s_axi_wdata   ( m31_axi_wdata   ),
  .s_axi_wstrb   ( m31_axi_wstrb   ),
  .s_axi_wlast   ( m31_axi_wlast   ),
  .s_axi_bvalid  ( m31_axi_bvalid  ),
  .s_axi_bready  ( m31_axi_bready  ),
  .s_axi_arvalid ( m31_axi_arvalid ),
  .s_axi_arready ( m31_axi_arready ),
  .s_axi_araddr  ( m31_axi_araddr  ),
  .s_axi_arlen   ( m31_axi_arlen   ),
  .s_axi_rvalid  ( m31_axi_rvalid  ),
  .s_axi_rready  ( m31_axi_rready  ),
  .s_axi_rdata   ( m31_axi_rdata   ),
  .s_axi_rlast   ( m31_axi_rlast   )
);


slv_m31_axi_vip_slv_mem_t   m31_axi;
slv_m31_axi_vip_slv_t   m31_axi_slv;

parameter NUM_AXIS_MST = 0;
parameter NUM_AXIS_SLV = 0;
parameter NUM_AXIS_PAIRS = 0;
bit               error_found = 0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m00_axi
bit [63:0] axi00_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m01_axi
bit [63:0] axi01_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m02_axi
bit [63:0] axi02_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m03_axi
bit [63:0] axi03_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m04_axi
bit [63:0] axi04_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m05_axi
bit [63:0] axi05_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m06_axi
bit [63:0] axi06_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m07_axi
bit [63:0] axi07_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m08_axi
bit [63:0] axi08_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m09_axi
bit [63:0] axi09_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m10_axi
bit [63:0] axi10_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m11_axi
bit [63:0] axi11_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m12_axi
bit [63:0] axi12_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m13_axi
bit [63:0] axi13_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m14_axi
bit [63:0] axi14_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m15_axi
bit [63:0] axi15_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m16_axi
bit [63:0] axi16_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m17_axi
bit [63:0] axi17_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m18_axi
bit [63:0] axi18_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m19_axi
bit [63:0] axi19_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m20_axi
bit [63:0] axi20_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m21_axi
bit [63:0] axi21_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m22_axi
bit [63:0] axi22_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m23_axi
bit [63:0] axi23_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m24_axi
bit [63:0] axi24_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m25_axi
bit [63:0] axi25_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m26_axi
bit [63:0] axi26_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m27_axi
bit [63:0] axi27_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m28_axi
bit [63:0] axi28_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m29_axi
bit [63:0] axi29_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m30_axi
bit [63:0] axi30_ptr0_ptr = 64'h0;

///////////////////////////////////////////////////////////////////////////
// Pointer for interface : m31_axi
bit [63:0] axi31_ptr0_ptr = 64'h0;

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m00_axi memory.
// write graph data
function void m00_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_0.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m00_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m01_axi memory.
function void m01_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_1.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m01_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m02_axi memory.
function void m02_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_2.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m02_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m03_axi memory.
function void m03_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_3.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m03_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m04_axi memory.
function void m04_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_4.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m04_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m05_axi memory.
function void m05_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_5.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m05_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m06_axi memory.
function void m06_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_6.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m06_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m07_axi memory.
function void m07_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_7.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m07_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m08_axi memory.
function void m08_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_8.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m08_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m09_axi memory.
function void m09_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_9.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m09_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m10_axi memory.
function void m10_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_10.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m10_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m11_axi memory.
function void m11_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_11.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m11_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m12_axi memory.
function void m12_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_12.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m12_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m13_axi memory.
function void m13_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_13.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m13_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m14_axi memory.
function void m14_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_14.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m14_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m15_axi memory.
function void m15_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_15.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m15_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m16_axi memory.
function void m16_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_16.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m16_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m17_axi memory.
function void m17_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_17.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m17_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m18_axi memory.
function void m18_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_18.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m18_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m19_axi memory.
function void m19_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_19.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m19_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m20_axi memory.
function void m20_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_20.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m20_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m21_axi memory.
function void m21_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_21.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m21_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m22_axi memory.
function void m22_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_22.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m22_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m23_axi memory.
function void m23_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_23.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m23_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m24_axi memory.
function void m24_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_24.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m24_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m25_axi memory.
function void m25_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_25.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m25_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m26_axi memory.
function void m26_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_26.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m26_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m27_axi memory.
function void m27_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_27.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m27_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m28_axi memory.
function void m28_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_28.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m28_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m29_axi memory.
function void m29_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_29.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m29_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m30_axi memory.
function void m30_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_30.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m30_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Backdoor fill the m31_axi memory.
function void m31_axi_fill_memory(
  input bit [63:0] ptr,
  input integer    length
);
  integer fd;
  reg [31 : 0] data;
  fd = $fopen({file_location,"edge_channel_small_31.txt"}, "r");
  if (!fd && length) begin
    $finish();
  end
  for (longint unsigned slot = 0; slot < length; slot++) begin
    $fscanf(fd, "%d", data);
    m31_axi.mem_model.backdoor_memory_write_4byte(ptr + (slot * 4), data);
  end
endfunction

task automatic system_reset_sequence(input integer unsigned width = 20);
  $display("%t : Starting System Reset Sequence", $time);
  fork
    ap_rst_n_sequence(25);
    
    
  join

endtask


/////////////////////////////////////////////////////////////////////////////////////////////////
// Generate a random 32bit number
function bit [31:0] get_random_4bytes();
  bit [31:0] rptr;
  ptr_random_failed: assert(std::randomize(rptr));
  return(rptr);
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Generate a random 64bit 4k aligned address pointer.
function bit [63:0] get_random_ptr();
  bit [63:0] rptr;
  ptr_random_failed: assert(std::randomize(rptr));
  rptr[31:0] &= ~(32'h00000fff);
  return(rptr);
endfunction

/////////////////////////////////////////////////////////////////////////////////////////////////
// Control interface non-blocking write
// The task will return when the transaction has been accepted by the driver. It will be some
// amount of time before it will appear on the interface.
task automatic write_register (input bit [31:0] addr_in, input bit [31:0] data);
  axi_transaction   wr_xfer;
  wr_xfer = ctrl.wr_driver.create_transaction("wr_xfer");
  assert(wr_xfer.randomize() with {addr == addr_in;});
  wr_xfer.set_data_beat(0, data);
  ctrl.wr_driver.send(wr_xfer);
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Control interface blocking write
// The task will return when the BRESP has been returned from the kernel.
task automatic blocking_write_register (input bit [31:0] addr_in, input bit [31:0] data);
  axi_transaction   wr_xfer;
  axi_transaction   wr_rsp;
  wr_xfer = ctrl.wr_driver.create_transaction("wr_xfer");
  wr_xfer.set_driver_return_item_policy(XIL_AXI_PAYLOAD_RETURN);
  assert(wr_xfer.randomize() with {addr == addr_in;});
  wr_xfer.set_data_beat(0, data);
  ctrl.wr_driver.send(wr_xfer);
  ctrl.wr_driver.wait_rsp(wr_rsp);
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Control interface blocking read
// The task will return when the BRESP has been returned from the kernel.
task automatic read_register (input bit [31:0] addr, output bit [31:0] rddata);
  axi_transaction   rd_xfer;
  axi_transaction   rd_rsp;
  bit [31:0] rd_value;
  rd_xfer = ctrl.rd_driver.create_transaction("rd_xfer");
  rd_xfer.set_addr(addr);
  rd_xfer.set_driver_return_item_policy(XIL_AXI_PAYLOAD_RETURN);
  ctrl.rd_driver.send(rd_xfer);
  ctrl.rd_driver.wait_rsp(rd_rsp);
  rd_value = rd_rsp.get_data_beat(0);
  rddata = rd_value;
endtask



/////////////////////////////////////////////////////////////////////////////////////////////////
// Poll the Control interface status register.
// This will poll until the DONE flag in the status register is asserted.
task automatic poll_done_register ();
  bit [31:0] rd_value;
  do begin
    read_register(KRNL_CTRL_REG_ADDR, rd_value);
  end while ((rd_value & CTRL_DONE_MASK) == 0);
endtask

// This will poll until the IDLE flag in the status register is asserted.
task automatic poll_idle_register ();
  bit [31:0] rd_value;
  do begin
    read_register(KRNL_CTRL_REG_ADDR, rd_value);
  end while ((rd_value & CTRL_IDLE_MASK) == 0);
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Write to the control registers to enable the triggering of interrupts for the kernel
task automatic enable_interrupts();
  $display("Starting: Enabling Interrupts....");
  write_register(KRNL_GIE_REG_ADDR, GIE_GIE_MASK);
  write_register(KRNL_IER_REG_ADDR, IER_DONE_MASK);
  $display("Finished: Interrupts enabled.");
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Disabled the interrupts.
task automatic disable_interrupts();
  $display("Starting: Disable Interrupts....");
  write_register(KRNL_GIE_REG_ADDR, 32'h0);
  write_register(KRNL_IER_REG_ADDR, 32'h0);
  $display("Finished: Interrupts disabled.");
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
//When the interrupt is asserted, read the correct registers and clear the asserted interrupt.
task automatic service_interrupts();
  bit [31:0] rd_value;
  $display("Starting Servicing interrupts....");
  read_register(KRNL_CTRL_REG_ADDR, rd_value);
  $display("Control Register: 0x%0x", rd_value);

  blocking_write_register(KRNL_CTRL_REG_ADDR, rd_value);

  if ((rd_value & CTRL_DONE_MASK) == 0) begin
    $error("%t : DONE bit not asserted. Register value: (0x%0x)", $time, rd_value);
  end
  read_register(KRNL_ISR_REG_ADDR, rd_value);
  $display("Interrupt Status Register: 0x%0x", rd_value);
  blocking_write_register(KRNL_ISR_REG_ADDR, rd_value);
  $display("Finished Servicing interrupts");
endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Start the control VIP, SLAVE memory models and AXI4-Stream.
task automatic start_vips();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Control Master: ctrl");
  ctrl = new("ctrl", acc_kernel_tb.inst_control_acc_kernel_vip.inst.IF);
  ctrl.start_master();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m00_axi");
  m00_axi = new("m00_axi", acc_kernel_tb.inst_slv_m00_axi_vip.inst.IF);
  m00_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m01_axi");
  m01_axi = new("m01_axi", acc_kernel_tb.inst_slv_m01_axi_vip.inst.IF);
  m01_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m02_axi");
  m02_axi = new("m02_axi", acc_kernel_tb.inst_slv_m02_axi_vip.inst.IF);
  m02_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m03_axi");
  m03_axi = new("m03_axi", acc_kernel_tb.inst_slv_m03_axi_vip.inst.IF);
  m03_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m04_axi");
  m04_axi = new("m04_axi", acc_kernel_tb.inst_slv_m04_axi_vip.inst.IF);
  m04_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m05_axi");
  m05_axi = new("m05_axi", acc_kernel_tb.inst_slv_m05_axi_vip.inst.IF);
  m05_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m06_axi");
  m06_axi = new("m06_axi", acc_kernel_tb.inst_slv_m06_axi_vip.inst.IF);
  m06_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m07_axi");
  m07_axi = new("m07_axi", acc_kernel_tb.inst_slv_m07_axi_vip.inst.IF);
  m07_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m08_axi");
  m08_axi = new("m08_axi", acc_kernel_tb.inst_slv_m08_axi_vip.inst.IF);
  m08_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m09_axi");
  m09_axi = new("m09_axi", acc_kernel_tb.inst_slv_m09_axi_vip.inst.IF);
  m09_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m10_axi");
  m10_axi = new("m10_axi", acc_kernel_tb.inst_slv_m10_axi_vip.inst.IF);
  m10_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m11_axi");
  m11_axi = new("m11_axi", acc_kernel_tb.inst_slv_m11_axi_vip.inst.IF);
  m11_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m12_axi");
  m12_axi = new("m12_axi", acc_kernel_tb.inst_slv_m12_axi_vip.inst.IF);
  m12_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m13_axi");
  m13_axi = new("m13_axi", acc_kernel_tb.inst_slv_m13_axi_vip.inst.IF);
  m13_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m14_axi");
  m14_axi = new("m14_axi", acc_kernel_tb.inst_slv_m14_axi_vip.inst.IF);
  m14_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m15_axi");
  m15_axi = new("m15_axi", acc_kernel_tb.inst_slv_m15_axi_vip.inst.IF);
  m15_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m16_axi");
  m16_axi = new("m16_axi", acc_kernel_tb.inst_slv_m16_axi_vip.inst.IF);
  m16_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m17_axi");
  m17_axi = new("m17_axi", acc_kernel_tb.inst_slv_m17_axi_vip.inst.IF);
  m17_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m18_axi");
  m18_axi = new("m18_axi", acc_kernel_tb.inst_slv_m18_axi_vip.inst.IF);
  m18_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m19_axi");
  m19_axi = new("m19_axi", acc_kernel_tb.inst_slv_m19_axi_vip.inst.IF);
  m19_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m20_axi");
  m20_axi = new("m20_axi", acc_kernel_tb.inst_slv_m20_axi_vip.inst.IF);
  m20_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m21_axi");
  m21_axi = new("m21_axi", acc_kernel_tb.inst_slv_m21_axi_vip.inst.IF);
  m21_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m22_axi");
  m22_axi = new("m22_axi", acc_kernel_tb.inst_slv_m22_axi_vip.inst.IF);
  m22_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m23_axi");
  m23_axi = new("m23_axi", acc_kernel_tb.inst_slv_m23_axi_vip.inst.IF);
  m23_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m24_axi");
  m24_axi = new("m24_axi", acc_kernel_tb.inst_slv_m24_axi_vip.inst.IF);
  m24_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m25_axi");
  m25_axi = new("m25_axi", acc_kernel_tb.inst_slv_m25_axi_vip.inst.IF);
  m25_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m26_axi");
  m26_axi = new("m26_axi", acc_kernel_tb.inst_slv_m26_axi_vip.inst.IF);
  m26_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m27_axi");
  m27_axi = new("m27_axi", acc_kernel_tb.inst_slv_m27_axi_vip.inst.IF);
  m27_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m28_axi");
  m28_axi = new("m28_axi", acc_kernel_tb.inst_slv_m28_axi_vip.inst.IF);
  m28_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m29_axi");
  m29_axi = new("m29_axi", acc_kernel_tb.inst_slv_m29_axi_vip.inst.IF);
  m29_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m30_axi");
  m30_axi = new("m30_axi", acc_kernel_tb.inst_slv_m30_axi_vip.inst.IF);
  m30_axi.start_slave();

  $display("///////////////////////////////////////////////////////////////////////////");
  $display("Starting Memory slave: m31_axi");
  m31_axi = new("m31_axi", acc_kernel_tb.inst_slv_m31_axi_vip.inst.IF);
  m31_axi.start_slave();

endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// For each of the connected slave interfaces, set the Slave to not de-assert WREADY at any time.
// This will show the fastest outbound bandwidth from the WRITE channel.
task automatic slv_no_backpressure_wready();
  axi_ready_gen     rgen;
  $display("%t - Applying slv_no_backpressure_wready", $time);

  rgen = new("m00_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m00_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m01_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m01_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m02_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m02_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m03_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m03_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m04_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m04_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m05_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m05_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m06_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m06_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m07_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m07_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m08_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m08_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m09_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m09_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m10_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m10_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m11_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m11_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m12_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m12_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m13_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m13_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m14_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m14_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m15_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m15_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m16_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m16_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m17_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m17_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m18_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m18_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m19_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m19_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m20_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m20_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m21_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m21_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m22_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m22_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m23_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m23_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m24_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m24_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m25_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m25_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m26_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m26_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m27_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m27_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m28_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m28_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m29_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m29_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m30_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m30_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m31_axi_no_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_NO_BACKPRESSURE);
  m31_axi.wr_driver.set_wready_gen(rgen);

endtask


/////////////////////////////////////////////////////////////////////////////////////////////////
// For each of the connected slave interfaces, apply a WREADY policy to introduce backpressure.
// Based on the simulation seed the order/shape of the WREADY per-channel will be different.
task automatic slv_random_backpressure_wready();
  axi_ready_gen     rgen;
  $display("%t - Applying slv_random_backpressure_wready", $time);

  rgen = new("m00_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m00_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m01_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m01_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m02_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m02_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m03_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m03_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m04_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m04_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m05_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m05_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m06_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m06_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m07_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m07_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m08_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m08_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m09_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m09_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m10_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m10_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m11_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m11_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m12_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m12_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m13_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m13_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m14_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m14_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m15_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m15_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m16_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m16_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m17_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m17_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m18_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m18_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m19_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m19_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m20_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m20_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m21_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m21_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m22_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m22_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m23_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m23_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m24_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m24_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m25_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m25_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m26_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m26_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m27_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m27_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m28_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m28_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m29_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m29_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m30_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m30_axi.wr_driver.set_wready_gen(rgen);

  rgen = new("m31_axi_random_backpressure_wready");
  rgen.set_ready_policy(XIL_AXI_READY_GEN_RANDOM);
  rgen.set_low_time_range(0,12);
  rgen.set_high_time_range(1,12);
  rgen.set_event_count_range(3,5);
  m31_axi.wr_driver.set_wready_gen(rgen);

endtask


/////////////////////////////////////////////////////////////////////////////////////////////////
// For each of the connected slave interfaces, force the memory model to not insert any inter-beat
// gaps on the READ channel.
task automatic slv_no_delay_rvalid();
  $display("%t - Applying slv_no_delay_rvalid", $time);

  m00_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m00_axi.mem_model.set_inter_beat_gap(0);

  m01_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m01_axi.mem_model.set_inter_beat_gap(0);

  m02_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m02_axi.mem_model.set_inter_beat_gap(0);

  m03_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m03_axi.mem_model.set_inter_beat_gap(0);

  m04_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m04_axi.mem_model.set_inter_beat_gap(0);

  m05_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m05_axi.mem_model.set_inter_beat_gap(0);

  m06_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m06_axi.mem_model.set_inter_beat_gap(0);

  m07_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m07_axi.mem_model.set_inter_beat_gap(0);

  m08_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m08_axi.mem_model.set_inter_beat_gap(0);

  m09_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m09_axi.mem_model.set_inter_beat_gap(0);

  m10_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m10_axi.mem_model.set_inter_beat_gap(0);

  m11_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m11_axi.mem_model.set_inter_beat_gap(0);

  m12_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m12_axi.mem_model.set_inter_beat_gap(0);

  m13_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m13_axi.mem_model.set_inter_beat_gap(0);

  m14_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m14_axi.mem_model.set_inter_beat_gap(0);

  m15_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m15_axi.mem_model.set_inter_beat_gap(0);

  m16_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m16_axi.mem_model.set_inter_beat_gap(0);

  m17_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m17_axi.mem_model.set_inter_beat_gap(0);

  m18_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m18_axi.mem_model.set_inter_beat_gap(0);

  m19_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m19_axi.mem_model.set_inter_beat_gap(0);

  m20_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m20_axi.mem_model.set_inter_beat_gap(0);

  m21_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m21_axi.mem_model.set_inter_beat_gap(0);

  m22_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m22_axi.mem_model.set_inter_beat_gap(0);

  m23_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m23_axi.mem_model.set_inter_beat_gap(0);

  m24_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m24_axi.mem_model.set_inter_beat_gap(0);

  m25_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m25_axi.mem_model.set_inter_beat_gap(0);

  m26_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m26_axi.mem_model.set_inter_beat_gap(0);

  m27_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m27_axi.mem_model.set_inter_beat_gap(0);

  m28_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m28_axi.mem_model.set_inter_beat_gap(0);

  m29_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m29_axi.mem_model.set_inter_beat_gap(0);

  m30_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m30_axi.mem_model.set_inter_beat_gap(0);

  m31_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_FIXED);
  m31_axi.mem_model.set_inter_beat_gap(0);

endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// For each of the connected slave interfaces, Allow the memory model to insert any inter-beat
// gaps on the READ channel.
task automatic slv_random_delay_rvalid();
  $display("%t - Applying slv_random_delay_rvalid", $time);

  m00_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m00_axi.mem_model.set_inter_beat_gap_range(0,10);

  m01_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m01_axi.mem_model.set_inter_beat_gap_range(0,10);

  m02_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m02_axi.mem_model.set_inter_beat_gap_range(0,10);

  m03_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m03_axi.mem_model.set_inter_beat_gap_range(0,10);

  m04_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m04_axi.mem_model.set_inter_beat_gap_range(0,10);

  m05_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m05_axi.mem_model.set_inter_beat_gap_range(0,10);

  m06_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m06_axi.mem_model.set_inter_beat_gap_range(0,10);

  m07_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m07_axi.mem_model.set_inter_beat_gap_range(0,10);

  m08_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m08_axi.mem_model.set_inter_beat_gap_range(0,10);

  m09_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m09_axi.mem_model.set_inter_beat_gap_range(0,10);

  m10_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m10_axi.mem_model.set_inter_beat_gap_range(0,10);

  m11_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m11_axi.mem_model.set_inter_beat_gap_range(0,10);

  m12_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m12_axi.mem_model.set_inter_beat_gap_range(0,10);

  m13_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m13_axi.mem_model.set_inter_beat_gap_range(0,10);

  m14_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m14_axi.mem_model.set_inter_beat_gap_range(0,10);

  m15_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m15_axi.mem_model.set_inter_beat_gap_range(0,10);

  m16_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m16_axi.mem_model.set_inter_beat_gap_range(0,10);

  m17_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m17_axi.mem_model.set_inter_beat_gap_range(0,10);

  m18_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m18_axi.mem_model.set_inter_beat_gap_range(0,10);

  m19_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m19_axi.mem_model.set_inter_beat_gap_range(0,10);

  m20_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m20_axi.mem_model.set_inter_beat_gap_range(0,10);

  m21_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m21_axi.mem_model.set_inter_beat_gap_range(0,10);

  m22_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m22_axi.mem_model.set_inter_beat_gap_range(0,10);

  m23_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m23_axi.mem_model.set_inter_beat_gap_range(0,10);

  m24_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m24_axi.mem_model.set_inter_beat_gap_range(0,10);

  m25_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m25_axi.mem_model.set_inter_beat_gap_range(0,10);

  m26_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m26_axi.mem_model.set_inter_beat_gap_range(0,10);

  m27_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m27_axi.mem_model.set_inter_beat_gap_range(0,10);

  m28_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m28_axi.mem_model.set_inter_beat_gap_range(0,10);

  m29_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m29_axi.mem_model.set_inter_beat_gap_range(0,10);

  m30_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m30_axi.mem_model.set_inter_beat_gap_range(0,10);

  m31_axi.mem_model.set_inter_beat_gap_delay_policy(XIL_AXI_MEMORY_DELAY_RANDOM);
  m31_axi.mem_model.set_inter_beat_gap_range(0,10);

endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
// Check to ensure, following reset the value of the register is 0.
// Check that only the width of the register bits can be written.
task automatic check_register_value(input bit [31:0] addr_in, input integer unsigned register_width, output bit error_found);
  bit [31:0] rddata;
  bit [31:0] mask_data;
  error_found = 0;
  if (register_width < 32) begin
    mask_data = (1 << register_width) - 1;
  end else begin
    mask_data = 32'hffffffff;
  end
  read_register(addr_in, rddata);
  if (rddata != 32'h0) begin
    $error("Initial value mismatch: A:0x%0x : Expected 0x%x -> Got 0x%x", addr_in, 0, rddata);
    error_found = 1;
  end
  blocking_write_register(addr_in, 32'hffffffff);
  read_register(addr_in, rddata);
  if (rddata != mask_data) begin
    $error("Initial value mismatch: A:0x%0x : Expected 0x%x -> Got 0x%x", addr_in, mask_data, rddata);
    error_found = 1;
  end
endtask


/////////////////////////////////////////////////////////////////////////////////////////////////
// For each of the scalar registers, check:
// * reset value
// * correct number bits set on a write
task automatic check_scalar_registers(output bit error_found);
  bit tmp_error_found = 0;
  error_found = 0;
  $display("%t : Checking post reset values of scalar registers", $time);

  ///////////////////////////////////////////////////////////////////////////
  //Check ID 0: root_id (0x010)
  check_register_value(32'h010, 32, tmp_error_found);
  error_found |= tmp_error_found;

endtask

task automatic set_scalar_registers();
  $display("%t : Setting Scalar Registers registers", $time);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 0: root_id (0x010) -> 32'hffffffff (scalar)
  // write_register(32'h010, 32'hffffffff);
  write_register(32'h010, 32'h00000001); // set root_id=1

endtask

task automatic check_pointer_registers(output bit error_found);
  bit tmp_error_found = 0;
  ///////////////////////////////////////////////////////////////////////////
  //Check the reset states of the pointer registers.
  $display("%t : Checking post reset values of pointer registers", $time);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 1: axi00_ptr0 (0x018)
  check_register_value(32'h018, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 1: axi00_ptr0 (0x01c)
  check_register_value(32'h01c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 2: axi01_ptr0 (0x024)
  check_register_value(32'h024, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 2: axi01_ptr0 (0x028)
  check_register_value(32'h028, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 3: axi02_ptr0 (0x030)
  check_register_value(32'h030, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 3: axi02_ptr0 (0x034)
  check_register_value(32'h034, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 4: axi03_ptr0 (0x03c)
  check_register_value(32'h03c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 4: axi03_ptr0 (0x040)
  check_register_value(32'h040, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 5: axi04_ptr0 (0x048)
  check_register_value(32'h048, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 5: axi04_ptr0 (0x04c)
  check_register_value(32'h04c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 6: axi05_ptr0 (0x054)
  check_register_value(32'h054, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 6: axi05_ptr0 (0x058)
  check_register_value(32'h058, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 7: axi06_ptr0 (0x060)
  check_register_value(32'h060, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 7: axi06_ptr0 (0x064)
  check_register_value(32'h064, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 8: axi07_ptr0 (0x06c)
  check_register_value(32'h06c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 8: axi07_ptr0 (0x070)
  check_register_value(32'h070, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 9: axi08_ptr0 (0x078)
  check_register_value(32'h078, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 9: axi08_ptr0 (0x07c)
  check_register_value(32'h07c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 10: axi09_ptr0 (0x084)
  check_register_value(32'h084, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 10: axi09_ptr0 (0x088)
  check_register_value(32'h088, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 11: axi10_ptr0 (0x090)
  check_register_value(32'h090, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 11: axi10_ptr0 (0x094)
  check_register_value(32'h094, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 12: axi11_ptr0 (0x09c)
  check_register_value(32'h09c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 12: axi11_ptr0 (0x0a0)
  check_register_value(32'h0a0, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 13: axi12_ptr0 (0x0a8)
  check_register_value(32'h0a8, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 13: axi12_ptr0 (0x0ac)
  check_register_value(32'h0ac, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 14: axi13_ptr0 (0x0b4)
  check_register_value(32'h0b4, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 14: axi13_ptr0 (0x0b8)
  check_register_value(32'h0b8, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 15: axi14_ptr0 (0x0c0)
  check_register_value(32'h0c0, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 15: axi14_ptr0 (0x0c4)
  check_register_value(32'h0c4, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 16: axi15_ptr0 (0x0cc)
  check_register_value(32'h0cc, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 16: axi15_ptr0 (0x0d0)
  check_register_value(32'h0d0, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 17: axi16_ptr0 (0x0d8)
  check_register_value(32'h0d8, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 17: axi16_ptr0 (0x0dc)
  check_register_value(32'h0dc, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 18: axi17_ptr0 (0x0e4)
  check_register_value(32'h0e4, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 18: axi17_ptr0 (0x0e8)
  check_register_value(32'h0e8, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 19: axi18_ptr0 (0x0f0)
  check_register_value(32'h0f0, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 19: axi18_ptr0 (0x0f4)
  check_register_value(32'h0f4, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 20: axi19_ptr0 (0x0fc)
  check_register_value(32'h0fc, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 20: axi19_ptr0 (0x100)
  check_register_value(32'h100, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 21: axi20_ptr0 (0x108)
  check_register_value(32'h108, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 21: axi20_ptr0 (0x10c)
  check_register_value(32'h10c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 22: axi21_ptr0 (0x114)
  check_register_value(32'h114, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 22: axi21_ptr0 (0x118)
  check_register_value(32'h118, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 23: axi22_ptr0 (0x120)
  check_register_value(32'h120, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 23: axi22_ptr0 (0x124)
  check_register_value(32'h124, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 24: axi23_ptr0 (0x12c)
  check_register_value(32'h12c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 24: axi23_ptr0 (0x130)
  check_register_value(32'h130, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 25: axi24_ptr0 (0x138)
  check_register_value(32'h138, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 25: axi24_ptr0 (0x13c)
  check_register_value(32'h13c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 26: axi25_ptr0 (0x144)
  check_register_value(32'h144, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 26: axi25_ptr0 (0x148)
  check_register_value(32'h148, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 27: axi26_ptr0 (0x150)
  check_register_value(32'h150, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 27: axi26_ptr0 (0x154)
  check_register_value(32'h154, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 28: axi27_ptr0 (0x15c)
  check_register_value(32'h15c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 28: axi27_ptr0 (0x160)
  check_register_value(32'h160, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 29: axi28_ptr0 (0x168)
  check_register_value(32'h168, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 29: axi28_ptr0 (0x16c)
  check_register_value(32'h16c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 30: axi29_ptr0 (0x174)
  check_register_value(32'h174, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 30: axi29_ptr0 (0x178)
  check_register_value(32'h178, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 31: axi30_ptr0 (0x180)
  check_register_value(32'h180, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 31: axi30_ptr0 (0x184)
  check_register_value(32'h184, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 32: axi31_ptr0 (0x18c)
  check_register_value(32'h18c, 32, tmp_error_found);
  error_found |= tmp_error_found;

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 32: axi31_ptr0 (0x190)
  check_register_value(32'h190, 32, tmp_error_found);
  error_found |= tmp_error_found;

endtask

task automatic set_memory_pointers();
  ///////////////////////////////////////////////////////////////////////////
  //Randomly generate memory pointers.
  axi00_ptr0_ptr = get_random_ptr();
  axi01_ptr0_ptr = get_random_ptr();
  axi02_ptr0_ptr = get_random_ptr();
  axi03_ptr0_ptr = get_random_ptr();
  axi04_ptr0_ptr = get_random_ptr();
  axi05_ptr0_ptr = get_random_ptr();
  axi06_ptr0_ptr = get_random_ptr();
  axi07_ptr0_ptr = get_random_ptr();
  axi08_ptr0_ptr = get_random_ptr();
  axi09_ptr0_ptr = get_random_ptr();
  axi10_ptr0_ptr = get_random_ptr();
  axi11_ptr0_ptr = get_random_ptr();
  axi12_ptr0_ptr = get_random_ptr();
  axi13_ptr0_ptr = get_random_ptr();
  axi14_ptr0_ptr = get_random_ptr();
  axi15_ptr0_ptr = get_random_ptr();
  axi16_ptr0_ptr = get_random_ptr();
  axi17_ptr0_ptr = get_random_ptr();
  axi18_ptr0_ptr = get_random_ptr();
  axi19_ptr0_ptr = get_random_ptr();
  axi20_ptr0_ptr = get_random_ptr();
  axi21_ptr0_ptr = get_random_ptr();
  axi22_ptr0_ptr = get_random_ptr();
  axi23_ptr0_ptr = get_random_ptr();
  axi24_ptr0_ptr = get_random_ptr();
  axi25_ptr0_ptr = get_random_ptr();
  axi26_ptr0_ptr = get_random_ptr();
  axi27_ptr0_ptr = get_random_ptr();
  axi28_ptr0_ptr = get_random_ptr();
  axi29_ptr0_ptr = get_random_ptr();
  axi30_ptr0_ptr = get_random_ptr();
  axi31_ptr0_ptr = get_random_ptr();

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 1: axi00_ptr0 (0x018) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h018, axi00_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 1: axi00_ptr0 (0x01c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h01c, axi00_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 2: axi01_ptr0 (0x024) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h024, axi01_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 2: axi01_ptr0 (0x028) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h028, axi01_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 3: axi02_ptr0 (0x030) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h030, axi02_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 3: axi02_ptr0 (0x034) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h034, axi02_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 4: axi03_ptr0 (0x03c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h03c, axi03_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 4: axi03_ptr0 (0x040) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h040, axi03_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 5: axi04_ptr0 (0x048) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h048, axi04_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 5: axi04_ptr0 (0x04c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h04c, axi04_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 6: axi05_ptr0 (0x054) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h054, axi05_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 6: axi05_ptr0 (0x058) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h058, axi05_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 7: axi06_ptr0 (0x060) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h060, axi06_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 7: axi06_ptr0 (0x064) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h064, axi06_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 8: axi07_ptr0 (0x06c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h06c, axi07_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 8: axi07_ptr0 (0x070) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h070, axi07_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 9: axi08_ptr0 (0x078) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h078, axi08_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 9: axi08_ptr0 (0x07c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h07c, axi08_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 10: axi09_ptr0 (0x084) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h084, axi09_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 10: axi09_ptr0 (0x088) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h088, axi09_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 11: axi10_ptr0 (0x090) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h090, axi10_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 11: axi10_ptr0 (0x094) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h094, axi10_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 12: axi11_ptr0 (0x09c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h09c, axi11_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 12: axi11_ptr0 (0x0a0) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0a0, axi11_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 13: axi12_ptr0 (0x0a8) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0a8, axi12_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 13: axi12_ptr0 (0x0ac) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0ac, axi12_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 14: axi13_ptr0 (0x0b4) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0b4, axi13_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 14: axi13_ptr0 (0x0b8) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0b8, axi13_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 15: axi14_ptr0 (0x0c0) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0c0, axi14_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 15: axi14_ptr0 (0x0c4) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0c4, axi14_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 16: axi15_ptr0 (0x0cc) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0cc, axi15_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 16: axi15_ptr0 (0x0d0) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0d0, axi15_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 17: axi16_ptr0 (0x0d8) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0d8, axi16_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 17: axi16_ptr0 (0x0dc) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0dc, axi16_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 18: axi17_ptr0 (0x0e4) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0e4, axi17_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 18: axi17_ptr0 (0x0e8) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0e8, axi17_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 19: axi18_ptr0 (0x0f0) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0f0, axi18_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 19: axi18_ptr0 (0x0f4) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h0f4, axi18_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 20: axi19_ptr0 (0x0fc) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h0fc, axi19_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 20: axi19_ptr0 (0x100) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h100, axi19_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 21: axi20_ptr0 (0x108) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h108, axi20_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 21: axi20_ptr0 (0x10c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h10c, axi20_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 22: axi21_ptr0 (0x114) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h114, axi21_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 22: axi21_ptr0 (0x118) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h118, axi21_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 23: axi22_ptr0 (0x120) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h120, axi22_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 23: axi22_ptr0 (0x124) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h124, axi22_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 24: axi23_ptr0 (0x12c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h12c, axi23_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 24: axi23_ptr0 (0x130) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h130, axi23_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 25: axi24_ptr0 (0x138) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h138, axi24_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 25: axi24_ptr0 (0x13c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h13c, axi24_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 26: axi25_ptr0 (0x144) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h144, axi25_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 26: axi25_ptr0 (0x148) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h148, axi25_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 27: axi26_ptr0 (0x150) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h150, axi26_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 27: axi26_ptr0 (0x154) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h154, axi26_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 28: axi27_ptr0 (0x15c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h15c, axi27_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 28: axi27_ptr0 (0x160) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h160, axi27_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 29: axi28_ptr0 (0x168) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h168, axi28_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 29: axi28_ptr0 (0x16c) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h16c, axi28_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 30: axi29_ptr0 (0x174) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h174, axi29_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 30: axi29_ptr0 (0x178) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h178, axi29_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 31: axi30_ptr0 (0x180) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h180, axi30_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 31: axi30_ptr0 (0x184) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h184, axi30_ptr0_ptr[63:32]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 32: axi31_ptr0 (0x18c) -> Randomized 4k aligned address (Global memory, lower 32 bits)
  write_register(32'h18c, axi31_ptr0_ptr[31:0]);

  ///////////////////////////////////////////////////////////////////////////
  //Write ID 32: axi31_ptr0 (0x190) -> Randomized 4k aligned address (Global memory, upper 32 bits)
  write_register(32'h190, axi31_ptr0_ptr[63:32]);

endtask

task automatic backdoor_fill_memories();

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m00_axi_fill_memory(axi00_ptr0_ptr, 275247);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m01_axi_fill_memory(axi01_ptr0_ptr, 281195);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m02_axi_fill_memory(axi02_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m03_axi_fill_memory(axi03_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m04_axi_fill_memory(axi04_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m05_axi_fill_memory(axi05_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m06_axi_fill_memory(axi06_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m07_axi_fill_memory(axi07_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m08_axi_fill_memory(axi08_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m09_axi_fill_memory(axi09_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m10_axi_fill_memory(axi10_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m11_axi_fill_memory(axi11_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m12_axi_fill_memory(axi12_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m13_axi_fill_memory(axi13_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m14_axi_fill_memory(axi14_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m15_axi_fill_memory(axi15_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m16_axi_fill_memory(axi16_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m17_axi_fill_memory(axi17_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m18_axi_fill_memory(axi18_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m19_axi_fill_memory(axi19_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m20_axi_fill_memory(axi20_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m21_axi_fill_memory(axi21_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m22_axi_fill_memory(axi22_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m23_axi_fill_memory(axi23_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m24_axi_fill_memory(axi24_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m25_axi_fill_memory(axi25_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m26_axi_fill_memory(axi26_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m27_axi_fill_memory(axi27_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m28_axi_fill_memory(axi28_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m29_axi_fill_memory(axi29_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m30_axi_fill_memory(axi30_ptr0_ptr, 0);

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Backdoor fill the memory with the content.
  m31_axi_fill_memory(axi31_ptr0_ptr, 0);

endtask

function automatic bit check_kernel_result();
  bit [31:0]        ret_rd_value = 32'h0;
  bit error_found = 0;
  integer error_counter;
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m00_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m00_axi.mem_model.backdoor_memory_read_4byte(axi00_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m00_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi00_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m00_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi00_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m00_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m01_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m01_axi.mem_model.backdoor_memory_read_4byte(axi01_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m01_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi01_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m01_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi01_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m01_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m02_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m02_axi.mem_model.backdoor_memory_read_4byte(axi02_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m02_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi02_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m02_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi02_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m02_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m03_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m03_axi.mem_model.backdoor_memory_read_4byte(axi03_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m03_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi03_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m03_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi03_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m03_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m04_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m04_axi.mem_model.backdoor_memory_read_4byte(axi04_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m04_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi04_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m04_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi04_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m04_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m05_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m05_axi.mem_model.backdoor_memory_read_4byte(axi05_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m05_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi05_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m05_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi05_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m05_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m06_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m06_axi.mem_model.backdoor_memory_read_4byte(axi06_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m06_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi06_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m06_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi06_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m06_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m07_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m07_axi.mem_model.backdoor_memory_read_4byte(axi07_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m07_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi07_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m07_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi07_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m07_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m08_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m08_axi.mem_model.backdoor_memory_read_4byte(axi08_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m08_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi08_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m08_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi08_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m08_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m09_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m09_axi.mem_model.backdoor_memory_read_4byte(axi09_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m09_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi09_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m09_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi09_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m09_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m10_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m10_axi.mem_model.backdoor_memory_read_4byte(axi10_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m10_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi10_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m10_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi10_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m10_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m11_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m11_axi.mem_model.backdoor_memory_read_4byte(axi11_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m11_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi11_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m11_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi11_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m11_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m12_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m12_axi.mem_model.backdoor_memory_read_4byte(axi12_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m12_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi12_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m12_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi12_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m12_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m13_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m13_axi.mem_model.backdoor_memory_read_4byte(axi13_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m13_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi13_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m13_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi13_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m13_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m14_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m14_axi.mem_model.backdoor_memory_read_4byte(axi14_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m14_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi14_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m14_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi14_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m14_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m15_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m15_axi.mem_model.backdoor_memory_read_4byte(axi15_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m15_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi15_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m15_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi15_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m15_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m16_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m16_axi.mem_model.backdoor_memory_read_4byte(axi16_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m16_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi16_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m16_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi16_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m16_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m17_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m17_axi.mem_model.backdoor_memory_read_4byte(axi17_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m17_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi17_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m17_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi17_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m17_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m18_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m18_axi.mem_model.backdoor_memory_read_4byte(axi18_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m18_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi18_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m18_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi18_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m18_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m19_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m19_axi.mem_model.backdoor_memory_read_4byte(axi19_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m19_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi19_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m19_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi19_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m19_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m20_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m20_axi.mem_model.backdoor_memory_read_4byte(axi20_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m20_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi20_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m20_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi20_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m20_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m21_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m21_axi.mem_model.backdoor_memory_read_4byte(axi21_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m21_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi21_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m21_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi21_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m21_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m22_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m22_axi.mem_model.backdoor_memory_read_4byte(axi22_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m22_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi22_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m22_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi22_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m22_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m23_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m23_axi.mem_model.backdoor_memory_read_4byte(axi23_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m23_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi23_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m23_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi23_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m23_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m24_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m24_axi.mem_model.backdoor_memory_read_4byte(axi24_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m24_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi24_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m24_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi24_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m24_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m25_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m25_axi.mem_model.backdoor_memory_read_4byte(axi25_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m25_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi25_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m25_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi25_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m25_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m26_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m26_axi.mem_model.backdoor_memory_read_4byte(axi26_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m26_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi26_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m26_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi26_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m26_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m27_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m27_axi.mem_model.backdoor_memory_read_4byte(axi27_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m27_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi27_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m27_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi27_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m27_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m28_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m28_axi.mem_model.backdoor_memory_read_4byte(axi28_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m28_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi28_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m28_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi28_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m28_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m29_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m29_axi.mem_model.backdoor_memory_read_4byte(axi29_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m29_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi29_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m29_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi29_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m29_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m30_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m30_axi.mem_model.backdoor_memory_read_4byte(axi30_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m30_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi30_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m30_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi30_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m30_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  /////////////////////////////////////////////////////////////////////////////////////////////////
  // Checking memory connected to m31_axi
  for (longint unsigned slot = 0; slot < LP_MAX_LENGTH; slot++) begin
    ret_rd_value = m31_axi.mem_model.backdoor_memory_read_4byte(axi31_ptr0_ptr + (slot * 4));
    if (slot < LP_MAX_TRANSFER_LENGTH) begin
      if (ret_rd_value != (slot + 1)) begin
        $error("Memory Mismatch: m31_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi31_ptr0_ptr + (slot * 4), slot + 1, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end else begin
      if (ret_rd_value != slot) begin
        $error("Memory Mismatch: m31_axi : @0x%x : Expected 0x%x -> Got 0x%x ", axi31_ptr0_ptr + (slot * 4), slot, ret_rd_value);
        error_found |= 1;
        error_counter++;
      end
    end
    if (error_counter > 5) begin
      $display("Too many errors found. Exiting check of m31_axi.");
      slot = LP_MAX_LENGTH;
    end
  end
  error_counter = 0;

  return(error_found);
endfunction

bit choose_pressure_type = 0;
bit axis_choose_pressure_type = 0;
bit [0-1:0] axis_tlast_received;

/////////////////////////////////////////////////////////////////////////////////////////////////
// Set up the kernel for operation and set the kernel START bit.
// The task will poll the DONE bit and check the results when complete.
task automatic multiple_iteration(input integer unsigned num_iterations, output bit error_found);
  error_found = 0;

  $display("Starting: multiple_iteration");
  for (integer unsigned iter = 0; iter < num_iterations; iter++) begin

    
    $display("Starting iteration: %d / %d", iter+1, num_iterations);
    RAND_WREADY_PRESSURE_FAILED: assert(std::randomize(choose_pressure_type));
    case(choose_pressure_type)
      0: slv_no_backpressure_wready();
      1: slv_random_backpressure_wready();
    endcase
    RAND_RVALID_PRESSURE_FAILED: assert(std::randomize(choose_pressure_type));
    case(choose_pressure_type)
      0: slv_no_delay_rvalid();
      1: slv_random_delay_rvalid();
    endcase

    set_scalar_registers();
    set_memory_pointers();
    backdoor_fill_memories();
    // Check that Kernel is IDLE before starting.
    poll_idle_register();
    ///////////////////////////////////////////////////////////////////////////
    //Start transfers
    blocking_write_register(KRNL_CTRL_REG_ADDR, CTRL_START_MASK);

    ctrl.wait_drivers_idle();
    ///////////////////////////////////////////////////////////////////////////
    //Wait for interrupt being asserted or poll done register
    @(posedge interrupt);

    ///////////////////////////////////////////////////////////////////////////
    // Service the interrupt
    service_interrupts();
    wait(interrupt == 0);

    ///////////////////////////////////////////////////////////////////////////
    error_found |= check_kernel_result()   ;

    $display("Finished iteration: %d / %d", iter+1, num_iterations);
  end
 endtask

/////////////////////////////////////////////////////////////////////////////////////////////////
//Instantiate AXI4 LITE VIP
initial begin : STIMULUS
  #200000;
  start_vips();
  check_scalar_registers(error_found);
  if (error_found == 1) begin
    $display( "Test Failed!");
    $finish();
  end

  check_pointer_registers(error_found);
  if (error_found == 1) begin
    $display( "Test Failed!");
    $finish();
  end

  enable_interrupts();

  multiple_iteration(1, error_found);
  if (error_found == 1) begin
    $display( "Test Failed!");
    $finish();
  end

  multiple_iteration(5, error_found);

  if (error_found == 1) begin
    $display( "Test Failed!");
    $finish();
  end else begin
    $display( "Test completed successfully");
  end
  $finish;
end

endmodule
`default_nettype wire